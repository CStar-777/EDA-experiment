//megafunction wizard: %Altera SOPC Builder%
//GENERATION: STANDARD
//VERSION: WM1.0


//Legal Notice: (C)2021 Altera Corporation. All rights reserved.  Your
//use of Altera Corporation's design tools, logic functions and other
//software and tools, and its AMPP partner logic functions, and any
//output files any of the foregoing (including device programming or
//simulation files), and any associated documentation or information are
//expressly subject to the terms and conditions of the Altera Program
//License Subscription Agreement or other applicable license agreement,
//including, without limitation, that your use is for the sole purpose
//of programming logic devices manufactured by Altera and sold by Altera
//or its authorized distributors.  Please refer to the applicable
//agreement for further details.

// synthesis translate_off
`timescale 1ns / 1ps
// synthesis translate_on

// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module button_pio_s1_arbitrator (
                                  // inputs:
                                   button_pio_s1_irq,
                                   button_pio_s1_readdata,
                                   clk,
                                   cpu_0_data_master_address_to_slave,
                                   cpu_0_data_master_byteenable,
                                   cpu_0_data_master_latency_counter,
                                   cpu_0_data_master_read,
                                   cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                   cpu_0_data_master_write,
                                   cpu_0_data_master_writedata,
                                   reset_n,

                                  // outputs:
                                   button_pio_s1_address,
                                   button_pio_s1_chipselect,
                                   button_pio_s1_irq_from_sa,
                                   button_pio_s1_readdata_from_sa,
                                   button_pio_s1_reset_n,
                                   button_pio_s1_write_n,
                                   button_pio_s1_writedata,
                                   cpu_0_data_master_granted_button_pio_s1,
                                   cpu_0_data_master_qualified_request_button_pio_s1,
                                   cpu_0_data_master_read_data_valid_button_pio_s1,
                                   cpu_0_data_master_requests_button_pio_s1,
                                   d1_button_pio_s1_end_xfer
                                )
;

  output  [  1: 0] button_pio_s1_address;
  output           button_pio_s1_chipselect;
  output           button_pio_s1_irq_from_sa;
  output  [  7: 0] button_pio_s1_readdata_from_sa;
  output           button_pio_s1_reset_n;
  output           button_pio_s1_write_n;
  output  [  7: 0] button_pio_s1_writedata;
  output           cpu_0_data_master_granted_button_pio_s1;
  output           cpu_0_data_master_qualified_request_button_pio_s1;
  output           cpu_0_data_master_read_data_valid_button_pio_s1;
  output           cpu_0_data_master_requests_button_pio_s1;
  output           d1_button_pio_s1_end_xfer;
  input            button_pio_s1_irq;
  input   [  7: 0] button_pio_s1_readdata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_allgrants;
  wire             button_pio_s1_allow_new_arb_cycle;
  wire             button_pio_s1_any_bursting_master_saved_grant;
  wire             button_pio_s1_any_continuerequest;
  wire             button_pio_s1_arb_counter_enable;
  reg     [  1: 0] button_pio_s1_arb_share_counter;
  wire    [  1: 0] button_pio_s1_arb_share_counter_next_value;
  wire    [  1: 0] button_pio_s1_arb_share_set_values;
  wire             button_pio_s1_beginbursttransfer_internal;
  wire             button_pio_s1_begins_xfer;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_end_xfer;
  wire             button_pio_s1_firsttransfer;
  wire             button_pio_s1_grant_vector;
  wire             button_pio_s1_in_a_read_cycle;
  wire             button_pio_s1_in_a_write_cycle;
  wire             button_pio_s1_irq_from_sa;
  wire             button_pio_s1_master_qreq_vector;
  wire             button_pio_s1_non_bursting_master_requests;
  wire             button_pio_s1_pretend_byte_enable;
  wire    [  7: 0] button_pio_s1_readdata_from_sa;
  reg              button_pio_s1_reg_firsttransfer;
  wire             button_pio_s1_reset_n;
  reg              button_pio_s1_slavearbiterlockenable;
  wire             button_pio_s1_slavearbiterlockenable2;
  wire             button_pio_s1_unreg_firsttransfer;
  wire             button_pio_s1_waits_for_read;
  wire             button_pio_s1_waits_for_write;
  wire             button_pio_s1_write_n;
  wire    [  7: 0] button_pio_s1_writedata;
  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_button_pio_s1;
  wire             cpu_0_data_master_qualified_request_button_pio_s1;
  wire             cpu_0_data_master_read_data_valid_button_pio_s1;
  wire             cpu_0_data_master_requests_button_pio_s1;
  wire             cpu_0_data_master_saved_grant_button_pio_s1;
  reg              d1_button_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_button_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 24: 0] shifted_address_to_button_pio_s1_from_cpu_0_data_master;
  wire             wait_for_button_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~button_pio_s1_end_xfer;
    end


  assign button_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_button_pio_s1));
  //assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_readdata_from_sa = button_pio_s1_readdata;

  assign cpu_0_data_master_requests_button_pio_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801050) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //button_pio_s1_arb_share_counter set values, which is an e_mux
  assign button_pio_s1_arb_share_set_values = 1;

  //button_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign button_pio_s1_non_bursting_master_requests = cpu_0_data_master_requests_button_pio_s1;

  //button_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign button_pio_s1_any_bursting_master_saved_grant = 0;

  //button_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign button_pio_s1_arb_share_counter_next_value = button_pio_s1_firsttransfer ? (button_pio_s1_arb_share_set_values - 1) : |button_pio_s1_arb_share_counter ? (button_pio_s1_arb_share_counter - 1) : 0;

  //button_pio_s1_allgrants all slave grants, which is an e_mux
  assign button_pio_s1_allgrants = |button_pio_s1_grant_vector;

  //button_pio_s1_end_xfer assignment, which is an e_assign
  assign button_pio_s1_end_xfer = ~(button_pio_s1_waits_for_read | button_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_button_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_button_pio_s1 = button_pio_s1_end_xfer & (~button_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //button_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign button_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_button_pio_s1 & button_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests);

  //button_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_arb_share_counter <= 0;
      else if (button_pio_s1_arb_counter_enable)
          button_pio_s1_arb_share_counter <= button_pio_s1_arb_share_counter_next_value;
    end


  //button_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_slavearbiterlockenable <= 0;
      else if ((|button_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_button_pio_s1) | (end_xfer_arb_share_counter_term_button_pio_s1 & ~button_pio_s1_non_bursting_master_requests))
          button_pio_s1_slavearbiterlockenable <= |button_pio_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master button_pio/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = button_pio_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //button_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign button_pio_s1_slavearbiterlockenable2 = |button_pio_s1_arb_share_counter_next_value;

  //cpu_0/data_master button_pio/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = button_pio_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //button_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign button_pio_s1_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_button_pio_s1 = cpu_0_data_master_requests_button_pio_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_button_pio_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_button_pio_s1 = cpu_0_data_master_granted_button_pio_s1 & cpu_0_data_master_read & ~button_pio_s1_waits_for_read;

  //button_pio_s1_writedata mux, which is an e_mux
  assign button_pio_s1_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_button_pio_s1 = cpu_0_data_master_qualified_request_button_pio_s1;

  //cpu_0/data_master saved-grant button_pio/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_button_pio_s1 = cpu_0_data_master_requests_button_pio_s1;

  //allow new arb cycle for button_pio/s1, which is an e_assign
  assign button_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign button_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign button_pio_s1_master_qreq_vector = 1;

  //button_pio_s1_reset_n assignment, which is an e_assign
  assign button_pio_s1_reset_n = reset_n;

  assign button_pio_s1_chipselect = cpu_0_data_master_granted_button_pio_s1;
  //button_pio_s1_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_firsttransfer = button_pio_s1_begins_xfer ? button_pio_s1_unreg_firsttransfer : button_pio_s1_reg_firsttransfer;

  //button_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign button_pio_s1_unreg_firsttransfer = ~(button_pio_s1_slavearbiterlockenable & button_pio_s1_any_continuerequest);

  //button_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          button_pio_s1_reg_firsttransfer <= 1'b1;
      else if (button_pio_s1_begins_xfer)
          button_pio_s1_reg_firsttransfer <= button_pio_s1_unreg_firsttransfer;
    end


  //button_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign button_pio_s1_beginbursttransfer_internal = button_pio_s1_begins_xfer;

  //~button_pio_s1_write_n assignment, which is an e_mux
  assign button_pio_s1_write_n = ~(((cpu_0_data_master_granted_button_pio_s1 & cpu_0_data_master_write)) & button_pio_s1_pretend_byte_enable);

  assign shifted_address_to_button_pio_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //button_pio_s1_address mux, which is an e_mux
  assign button_pio_s1_address = shifted_address_to_button_pio_s1_from_cpu_0_data_master >> 2;

  //d1_button_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_button_pio_s1_end_xfer <= 1;
      else 
        d1_button_pio_s1_end_xfer <= button_pio_s1_end_xfer;
    end


  //button_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_read = button_pio_s1_in_a_read_cycle & button_pio_s1_begins_xfer;

  //button_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_read_cycle = cpu_0_data_master_granted_button_pio_s1 & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = button_pio_s1_in_a_read_cycle;

  //button_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign button_pio_s1_waits_for_write = button_pio_s1_in_a_write_cycle & 0;

  //button_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign button_pio_s1_in_a_write_cycle = cpu_0_data_master_granted_button_pio_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = button_pio_s1_in_a_write_cycle;

  assign wait_for_button_pio_s1_counter = 0;
  //button_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  assign button_pio_s1_pretend_byte_enable = (cpu_0_data_master_granted_button_pio_s1)? cpu_0_data_master_byteenable :
    -1;

  //assign button_pio_s1_irq_from_sa = button_pio_s1_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign button_pio_s1_irq_from_sa = button_pio_s1_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //button_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module col_s1_arbitrator (
                           // inputs:
                            clk,
                            col_s1_readdata,
                            cpu_0_data_master_address_to_slave,
                            cpu_0_data_master_latency_counter,
                            cpu_0_data_master_read,
                            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                            cpu_0_data_master_write,
                            cpu_0_data_master_writedata,
                            reset_n,

                           // outputs:
                            col_s1_address,
                            col_s1_chipselect,
                            col_s1_readdata_from_sa,
                            col_s1_reset_n,
                            col_s1_write_n,
                            col_s1_writedata,
                            cpu_0_data_master_granted_col_s1,
                            cpu_0_data_master_qualified_request_col_s1,
                            cpu_0_data_master_read_data_valid_col_s1,
                            cpu_0_data_master_requests_col_s1,
                            d1_col_s1_end_xfer
                         )
;

  output  [  1: 0] col_s1_address;
  output           col_s1_chipselect;
  output  [  3: 0] col_s1_readdata_from_sa;
  output           col_s1_reset_n;
  output           col_s1_write_n;
  output  [  3: 0] col_s1_writedata;
  output           cpu_0_data_master_granted_col_s1;
  output           cpu_0_data_master_qualified_request_col_s1;
  output           cpu_0_data_master_read_data_valid_col_s1;
  output           cpu_0_data_master_requests_col_s1;
  output           d1_col_s1_end_xfer;
  input            clk;
  input   [  3: 0] col_s1_readdata;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input            reset_n;

  wire    [  1: 0] col_s1_address;
  wire             col_s1_allgrants;
  wire             col_s1_allow_new_arb_cycle;
  wire             col_s1_any_bursting_master_saved_grant;
  wire             col_s1_any_continuerequest;
  wire             col_s1_arb_counter_enable;
  reg     [  1: 0] col_s1_arb_share_counter;
  wire    [  1: 0] col_s1_arb_share_counter_next_value;
  wire    [  1: 0] col_s1_arb_share_set_values;
  wire             col_s1_beginbursttransfer_internal;
  wire             col_s1_begins_xfer;
  wire             col_s1_chipselect;
  wire             col_s1_end_xfer;
  wire             col_s1_firsttransfer;
  wire             col_s1_grant_vector;
  wire             col_s1_in_a_read_cycle;
  wire             col_s1_in_a_write_cycle;
  wire             col_s1_master_qreq_vector;
  wire             col_s1_non_bursting_master_requests;
  wire    [  3: 0] col_s1_readdata_from_sa;
  reg              col_s1_reg_firsttransfer;
  wire             col_s1_reset_n;
  reg              col_s1_slavearbiterlockenable;
  wire             col_s1_slavearbiterlockenable2;
  wire             col_s1_unreg_firsttransfer;
  wire             col_s1_waits_for_read;
  wire             col_s1_waits_for_write;
  wire             col_s1_write_n;
  wire    [  3: 0] col_s1_writedata;
  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_col_s1;
  wire             cpu_0_data_master_qualified_request_col_s1;
  wire             cpu_0_data_master_read_data_valid_col_s1;
  wire             cpu_0_data_master_requests_col_s1;
  wire             cpu_0_data_master_saved_grant_col_s1;
  reg              d1_col_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_col_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [ 24: 0] shifted_address_to_col_s1_from_cpu_0_data_master;
  wire             wait_for_col_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~col_s1_end_xfer;
    end


  assign col_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_col_s1));
  //assign col_s1_readdata_from_sa = col_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign col_s1_readdata_from_sa = col_s1_readdata;

  assign cpu_0_data_master_requests_col_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010c0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //col_s1_arb_share_counter set values, which is an e_mux
  assign col_s1_arb_share_set_values = 1;

  //col_s1_non_bursting_master_requests mux, which is an e_mux
  assign col_s1_non_bursting_master_requests = cpu_0_data_master_requests_col_s1;

  //col_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign col_s1_any_bursting_master_saved_grant = 0;

  //col_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign col_s1_arb_share_counter_next_value = col_s1_firsttransfer ? (col_s1_arb_share_set_values - 1) : |col_s1_arb_share_counter ? (col_s1_arb_share_counter - 1) : 0;

  //col_s1_allgrants all slave grants, which is an e_mux
  assign col_s1_allgrants = |col_s1_grant_vector;

  //col_s1_end_xfer assignment, which is an e_assign
  assign col_s1_end_xfer = ~(col_s1_waits_for_read | col_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_col_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_col_s1 = col_s1_end_xfer & (~col_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //col_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign col_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_col_s1 & col_s1_allgrants) | (end_xfer_arb_share_counter_term_col_s1 & ~col_s1_non_bursting_master_requests);

  //col_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          col_s1_arb_share_counter <= 0;
      else if (col_s1_arb_counter_enable)
          col_s1_arb_share_counter <= col_s1_arb_share_counter_next_value;
    end


  //col_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          col_s1_slavearbiterlockenable <= 0;
      else if ((|col_s1_master_qreq_vector & end_xfer_arb_share_counter_term_col_s1) | (end_xfer_arb_share_counter_term_col_s1 & ~col_s1_non_bursting_master_requests))
          col_s1_slavearbiterlockenable <= |col_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master col/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = col_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //col_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign col_s1_slavearbiterlockenable2 = |col_s1_arb_share_counter_next_value;

  //cpu_0/data_master col/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = col_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //col_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign col_s1_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_col_s1 = cpu_0_data_master_requests_col_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_col_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_col_s1 = cpu_0_data_master_granted_col_s1 & cpu_0_data_master_read & ~col_s1_waits_for_read;

  //col_s1_writedata mux, which is an e_mux
  assign col_s1_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_col_s1 = cpu_0_data_master_qualified_request_col_s1;

  //cpu_0/data_master saved-grant col/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_col_s1 = cpu_0_data_master_requests_col_s1;

  //allow new arb cycle for col/s1, which is an e_assign
  assign col_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign col_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign col_s1_master_qreq_vector = 1;

  //col_s1_reset_n assignment, which is an e_assign
  assign col_s1_reset_n = reset_n;

  assign col_s1_chipselect = cpu_0_data_master_granted_col_s1;
  //col_s1_firsttransfer first transaction, which is an e_assign
  assign col_s1_firsttransfer = col_s1_begins_xfer ? col_s1_unreg_firsttransfer : col_s1_reg_firsttransfer;

  //col_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign col_s1_unreg_firsttransfer = ~(col_s1_slavearbiterlockenable & col_s1_any_continuerequest);

  //col_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          col_s1_reg_firsttransfer <= 1'b1;
      else if (col_s1_begins_xfer)
          col_s1_reg_firsttransfer <= col_s1_unreg_firsttransfer;
    end


  //col_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign col_s1_beginbursttransfer_internal = col_s1_begins_xfer;

  //~col_s1_write_n assignment, which is an e_mux
  assign col_s1_write_n = ~(cpu_0_data_master_granted_col_s1 & cpu_0_data_master_write);

  assign shifted_address_to_col_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //col_s1_address mux, which is an e_mux
  assign col_s1_address = shifted_address_to_col_s1_from_cpu_0_data_master >> 2;

  //d1_col_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_col_s1_end_xfer <= 1;
      else 
        d1_col_s1_end_xfer <= col_s1_end_xfer;
    end


  //col_s1_waits_for_read in a cycle, which is an e_mux
  assign col_s1_waits_for_read = col_s1_in_a_read_cycle & col_s1_begins_xfer;

  //col_s1_in_a_read_cycle assignment, which is an e_assign
  assign col_s1_in_a_read_cycle = cpu_0_data_master_granted_col_s1 & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = col_s1_in_a_read_cycle;

  //col_s1_waits_for_write in a cycle, which is an e_mux
  assign col_s1_waits_for_write = col_s1_in_a_write_cycle & 0;

  //col_s1_in_a_write_cycle assignment, which is an e_assign
  assign col_s1_in_a_write_cycle = cpu_0_data_master_granted_col_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = col_s1_in_a_write_cycle;

  assign wait_for_col_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //col/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_jtag_debug_module_arbitrator (
                                            // inputs:
                                             clk,
                                             cpu_0_data_master_address_to_slave,
                                             cpu_0_data_master_byteenable,
                                             cpu_0_data_master_debugaccess,
                                             cpu_0_data_master_latency_counter,
                                             cpu_0_data_master_read,
                                             cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                             cpu_0_data_master_write,
                                             cpu_0_data_master_writedata,
                                             cpu_0_instruction_master_address_to_slave,
                                             cpu_0_instruction_master_latency_counter,
                                             cpu_0_instruction_master_read,
                                             cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                             cpu_0_jtag_debug_module_readdata,
                                             cpu_0_jtag_debug_module_resetrequest,
                                             reset_n,

                                            // outputs:
                                             cpu_0_data_master_granted_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
                                             cpu_0_data_master_requests_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
                                             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
                                             cpu_0_jtag_debug_module_address,
                                             cpu_0_jtag_debug_module_begintransfer,
                                             cpu_0_jtag_debug_module_byteenable,
                                             cpu_0_jtag_debug_module_chipselect,
                                             cpu_0_jtag_debug_module_debugaccess,
                                             cpu_0_jtag_debug_module_readdata_from_sa,
                                             cpu_0_jtag_debug_module_reset,
                                             cpu_0_jtag_debug_module_reset_n,
                                             cpu_0_jtag_debug_module_resetrequest_from_sa,
                                             cpu_0_jtag_debug_module_write,
                                             cpu_0_jtag_debug_module_writedata,
                                             d1_cpu_0_jtag_debug_module_end_xfer
                                          )
;

  output           cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  output           cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  output           cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  output  [  8: 0] cpu_0_jtag_debug_module_address;
  output           cpu_0_jtag_debug_module_begintransfer;
  output  [  3: 0] cpu_0_jtag_debug_module_byteenable;
  output           cpu_0_jtag_debug_module_chipselect;
  output           cpu_0_jtag_debug_module_debugaccess;
  output  [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  output           cpu_0_jtag_debug_module_reset;
  output           cpu_0_jtag_debug_module_reset_n;
  output           cpu_0_jtag_debug_module_resetrequest_from_sa;
  output           cpu_0_jtag_debug_module_write;
  output  [ 31: 0] cpu_0_jtag_debug_module_writedata;
  output           d1_cpu_0_jtag_debug_module_end_xfer;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input            cpu_0_data_master_debugaccess;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata;
  input            cpu_0_jtag_debug_module_resetrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module;
  wire    [  8: 0] cpu_0_jtag_debug_module_address;
  wire             cpu_0_jtag_debug_module_allgrants;
  wire             cpu_0_jtag_debug_module_allow_new_arb_cycle;
  wire             cpu_0_jtag_debug_module_any_bursting_master_saved_grant;
  wire             cpu_0_jtag_debug_module_any_continuerequest;
  reg     [  1: 0] cpu_0_jtag_debug_module_arb_addend;
  wire             cpu_0_jtag_debug_module_arb_counter_enable;
  reg     [  1: 0] cpu_0_jtag_debug_module_arb_share_counter;
  wire    [  1: 0] cpu_0_jtag_debug_module_arb_share_counter_next_value;
  wire    [  1: 0] cpu_0_jtag_debug_module_arb_share_set_values;
  wire    [  1: 0] cpu_0_jtag_debug_module_arb_winner;
  wire             cpu_0_jtag_debug_module_arbitration_holdoff_internal;
  wire             cpu_0_jtag_debug_module_beginbursttransfer_internal;
  wire             cpu_0_jtag_debug_module_begins_xfer;
  wire             cpu_0_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_0_jtag_debug_module_byteenable;
  wire             cpu_0_jtag_debug_module_chipselect;
  wire    [  3: 0] cpu_0_jtag_debug_module_chosen_master_double_vector;
  wire    [  1: 0] cpu_0_jtag_debug_module_chosen_master_rot_left;
  wire             cpu_0_jtag_debug_module_debugaccess;
  wire             cpu_0_jtag_debug_module_end_xfer;
  wire             cpu_0_jtag_debug_module_firsttransfer;
  wire    [  1: 0] cpu_0_jtag_debug_module_grant_vector;
  wire             cpu_0_jtag_debug_module_in_a_read_cycle;
  wire             cpu_0_jtag_debug_module_in_a_write_cycle;
  wire    [  1: 0] cpu_0_jtag_debug_module_master_qreq_vector;
  wire             cpu_0_jtag_debug_module_non_bursting_master_requests;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  reg              cpu_0_jtag_debug_module_reg_firsttransfer;
  wire             cpu_0_jtag_debug_module_reset;
  wire             cpu_0_jtag_debug_module_reset_n;
  wire             cpu_0_jtag_debug_module_resetrequest_from_sa;
  reg     [  1: 0] cpu_0_jtag_debug_module_saved_chosen_master_vector;
  reg              cpu_0_jtag_debug_module_slavearbiterlockenable;
  wire             cpu_0_jtag_debug_module_slavearbiterlockenable2;
  wire             cpu_0_jtag_debug_module_unreg_firsttransfer;
  wire             cpu_0_jtag_debug_module_waits_for_read;
  wire             cpu_0_jtag_debug_module_waits_for_write;
  wire             cpu_0_jtag_debug_module_write;
  wire    [ 31: 0] cpu_0_jtag_debug_module_writedata;
  reg              d1_cpu_0_jtag_debug_module_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module;
  wire    [ 24: 0] shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master;
  wire             wait_for_cpu_0_jtag_debug_module_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~cpu_0_jtag_debug_module_end_xfer;
    end


  assign cpu_0_jtag_debug_module_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module));
  //assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_jtag_debug_module_readdata_from_sa = cpu_0_jtag_debug_module_readdata;

  assign cpu_0_data_master_requests_cpu_0_jtag_debug_module = ({cpu_0_data_master_address_to_slave[24 : 11] , 11'b0} == 25'h1800800) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //cpu_0_jtag_debug_module_arb_share_counter set values, which is an e_mux
  assign cpu_0_jtag_debug_module_arb_share_set_values = 1;

  //cpu_0_jtag_debug_module_non_bursting_master_requests mux, which is an e_mux
  assign cpu_0_jtag_debug_module_non_bursting_master_requests = cpu_0_data_master_requests_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_requests_cpu_0_jtag_debug_module |
    cpu_0_data_master_requests_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0_jtag_debug_module_any_bursting_master_saved_grant mux, which is an e_mux
  assign cpu_0_jtag_debug_module_any_bursting_master_saved_grant = 0;

  //cpu_0_jtag_debug_module_arb_share_counter_next_value assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_arb_share_counter_next_value = cpu_0_jtag_debug_module_firsttransfer ? (cpu_0_jtag_debug_module_arb_share_set_values - 1) : |cpu_0_jtag_debug_module_arb_share_counter ? (cpu_0_jtag_debug_module_arb_share_counter - 1) : 0;

  //cpu_0_jtag_debug_module_allgrants all slave grants, which is an e_mux
  assign cpu_0_jtag_debug_module_allgrants = (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector) |
    (|cpu_0_jtag_debug_module_grant_vector);

  //cpu_0_jtag_debug_module_end_xfer assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_end_xfer = ~(cpu_0_jtag_debug_module_waits_for_read | cpu_0_jtag_debug_module_waits_for_write);

  //end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_end_xfer & (~cpu_0_jtag_debug_module_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //cpu_0_jtag_debug_module_arb_share_counter arbitration counter enable, which is an e_assign
  assign cpu_0_jtag_debug_module_arb_counter_enable = (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & cpu_0_jtag_debug_module_allgrants) | (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & ~cpu_0_jtag_debug_module_non_bursting_master_requests);

  //cpu_0_jtag_debug_module_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_arb_share_counter <= 0;
      else if (cpu_0_jtag_debug_module_arb_counter_enable)
          cpu_0_jtag_debug_module_arb_share_counter <= cpu_0_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_0_jtag_debug_module_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_slavearbiterlockenable <= 0;
      else if ((|cpu_0_jtag_debug_module_master_qreq_vector & end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module) | (end_xfer_arb_share_counter_term_cpu_0_jtag_debug_module & ~cpu_0_jtag_debug_module_non_bursting_master_requests))
          cpu_0_jtag_debug_module_slavearbiterlockenable <= |cpu_0_jtag_debug_module_arb_share_counter_next_value;
    end


  //cpu_0/data_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //cpu_0_jtag_debug_module_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign cpu_0_jtag_debug_module_slavearbiterlockenable2 = |cpu_0_jtag_debug_module_arb_share_counter_next_value;

  //cpu_0/data_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = cpu_0_jtag_debug_module_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master cpu_0/jtag_debug_module arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = cpu_0_jtag_debug_module_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted cpu_0/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module <= cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module ? 1 : (cpu_0_jtag_debug_module_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_cpu_0_jtag_debug_module & cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0_jtag_debug_module_any_continuerequest at least one master continues requesting, which is an e_mux
  assign cpu_0_jtag_debug_module_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module = cpu_0_data_master_requests_cpu_0_jtag_debug_module & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  assign cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_read & ~cpu_0_jtag_debug_module_waits_for_read;

  //cpu_0_jtag_debug_module_writedata mux, which is an e_mux
  assign cpu_0_jtag_debug_module_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_cpu_0_jtag_debug_module = (({cpu_0_instruction_master_address_to_slave[24 : 11] , 11'b0} == 25'h1800800) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted cpu_0/jtag_debug_module last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module <= cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module ? 1 : (cpu_0_jtag_debug_module_arbitration_holdoff_internal | ~cpu_0_data_master_requests_cpu_0_jtag_debug_module) ? 0 : last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_cpu_0_jtag_debug_module & cpu_0_data_master_requests_cpu_0_jtag_debug_module;

  assign cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module = cpu_0_instruction_master_requests_cpu_0_jtag_debug_module & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module = cpu_0_instruction_master_granted_cpu_0_jtag_debug_module & cpu_0_instruction_master_read & ~cpu_0_jtag_debug_module_waits_for_read;

  //allow new arb cycle for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;

  //cpu_0/instruction_master grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_instruction_master_granted_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_grant_vector[0];

  //cpu_0/instruction_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_arb_winner[0] && cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;

  //cpu_0/data_master assignment into master qualified-requests vector for cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_jtag_debug_module_master_qreq_vector[1] = cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;

  //cpu_0/data_master grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_data_master_granted_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_grant_vector[1];

  //cpu_0/data_master saved-grant cpu_0/jtag_debug_module, which is an e_assign
  assign cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module = cpu_0_jtag_debug_module_arb_winner[1] && cpu_0_data_master_requests_cpu_0_jtag_debug_module;

  //cpu_0/jtag_debug_module chosen-master double-vector, which is an e_assign
  assign cpu_0_jtag_debug_module_chosen_master_double_vector = {cpu_0_jtag_debug_module_master_qreq_vector, cpu_0_jtag_debug_module_master_qreq_vector} & ({~cpu_0_jtag_debug_module_master_qreq_vector, ~cpu_0_jtag_debug_module_master_qreq_vector} + cpu_0_jtag_debug_module_arb_addend);

  //stable onehot encoding of arb winner
  assign cpu_0_jtag_debug_module_arb_winner = (cpu_0_jtag_debug_module_allow_new_arb_cycle & | cpu_0_jtag_debug_module_grant_vector) ? cpu_0_jtag_debug_module_grant_vector : cpu_0_jtag_debug_module_saved_chosen_master_vector;

  //saved cpu_0_jtag_debug_module_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_saved_chosen_master_vector <= 0;
      else if (cpu_0_jtag_debug_module_allow_new_arb_cycle)
          cpu_0_jtag_debug_module_saved_chosen_master_vector <= |cpu_0_jtag_debug_module_grant_vector ? cpu_0_jtag_debug_module_grant_vector : cpu_0_jtag_debug_module_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign cpu_0_jtag_debug_module_grant_vector = {(cpu_0_jtag_debug_module_chosen_master_double_vector[1] | cpu_0_jtag_debug_module_chosen_master_double_vector[3]),
    (cpu_0_jtag_debug_module_chosen_master_double_vector[0] | cpu_0_jtag_debug_module_chosen_master_double_vector[2])};

  //cpu_0/jtag_debug_module chosen master rotated left, which is an e_assign
  assign cpu_0_jtag_debug_module_chosen_master_rot_left = (cpu_0_jtag_debug_module_arb_winner << 1) ? (cpu_0_jtag_debug_module_arb_winner << 1) : 1;

  //cpu_0/jtag_debug_module's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_arb_addend <= 1;
      else if (|cpu_0_jtag_debug_module_grant_vector)
          cpu_0_jtag_debug_module_arb_addend <= cpu_0_jtag_debug_module_end_xfer? cpu_0_jtag_debug_module_chosen_master_rot_left : cpu_0_jtag_debug_module_grant_vector;
    end


  assign cpu_0_jtag_debug_module_begintransfer = cpu_0_jtag_debug_module_begins_xfer;
  //assign lhs ~cpu_0_jtag_debug_module_reset of type reset_n to cpu_0_jtag_debug_module_reset_n, which is an e_assign
  assign cpu_0_jtag_debug_module_reset = ~cpu_0_jtag_debug_module_reset_n;

  //cpu_0_jtag_debug_module_reset_n assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_reset_n = reset_n;

  //assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign cpu_0_jtag_debug_module_resetrequest_from_sa = cpu_0_jtag_debug_module_resetrequest;

  assign cpu_0_jtag_debug_module_chipselect = cpu_0_data_master_granted_cpu_0_jtag_debug_module | cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  //cpu_0_jtag_debug_module_firsttransfer first transaction, which is an e_assign
  assign cpu_0_jtag_debug_module_firsttransfer = cpu_0_jtag_debug_module_begins_xfer ? cpu_0_jtag_debug_module_unreg_firsttransfer : cpu_0_jtag_debug_module_reg_firsttransfer;

  //cpu_0_jtag_debug_module_unreg_firsttransfer first transaction, which is an e_assign
  assign cpu_0_jtag_debug_module_unreg_firsttransfer = ~(cpu_0_jtag_debug_module_slavearbiterlockenable & cpu_0_jtag_debug_module_any_continuerequest);

  //cpu_0_jtag_debug_module_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_jtag_debug_module_reg_firsttransfer <= 1'b1;
      else if (cpu_0_jtag_debug_module_begins_xfer)
          cpu_0_jtag_debug_module_reg_firsttransfer <= cpu_0_jtag_debug_module_unreg_firsttransfer;
    end


  //cpu_0_jtag_debug_module_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign cpu_0_jtag_debug_module_beginbursttransfer_internal = cpu_0_jtag_debug_module_begins_xfer;

  //cpu_0_jtag_debug_module_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign cpu_0_jtag_debug_module_arbitration_holdoff_internal = cpu_0_jtag_debug_module_begins_xfer & cpu_0_jtag_debug_module_firsttransfer;

  //cpu_0_jtag_debug_module_write assignment, which is an e_mux
  assign cpu_0_jtag_debug_module_write = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_write;

  assign shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //cpu_0_jtag_debug_module_address mux, which is an e_mux
  assign cpu_0_jtag_debug_module_address = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? (shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_data_master >> 2) :
    (shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_cpu_0_jtag_debug_module_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_cpu_0_jtag_debug_module_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_cpu_0_jtag_debug_module_end_xfer <= 1;
      else 
        d1_cpu_0_jtag_debug_module_end_xfer <= cpu_0_jtag_debug_module_end_xfer;
    end


  //cpu_0_jtag_debug_module_waits_for_read in a cycle, which is an e_mux
  assign cpu_0_jtag_debug_module_waits_for_read = cpu_0_jtag_debug_module_in_a_read_cycle & cpu_0_jtag_debug_module_begins_xfer;

  //cpu_0_jtag_debug_module_in_a_read_cycle assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_in_a_read_cycle = (cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cpu_0_jtag_debug_module_in_a_read_cycle;

  //cpu_0_jtag_debug_module_waits_for_write in a cycle, which is an e_mux
  assign cpu_0_jtag_debug_module_waits_for_write = cpu_0_jtag_debug_module_in_a_write_cycle & 0;

  //cpu_0_jtag_debug_module_in_a_write_cycle assignment, which is an e_assign
  assign cpu_0_jtag_debug_module_in_a_write_cycle = cpu_0_data_master_granted_cpu_0_jtag_debug_module & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cpu_0_jtag_debug_module_in_a_write_cycle;

  assign wait_for_cpu_0_jtag_debug_module_counter = 0;
  //cpu_0_jtag_debug_module_byteenable byte enable port mux, which is an e_mux
  assign cpu_0_jtag_debug_module_byteenable = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? cpu_0_data_master_byteenable :
    -1;

  //debugaccess mux, which is an e_mux
  assign cpu_0_jtag_debug_module_debugaccess = (cpu_0_data_master_granted_cpu_0_jtag_debug_module)? cpu_0_data_master_debugaccess :
    0;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0/jtag_debug_module enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_cpu_0_jtag_debug_module + cpu_0_instruction_master_granted_cpu_0_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_cpu_0_jtag_debug_module + cpu_0_instruction_master_saved_grant_cpu_0_jtag_debug_module > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_data_master_arbitrator (
                                      // inputs:
                                       button_pio_s1_irq_from_sa,
                                       button_pio_s1_readdata_from_sa,
                                       cfi_flash_0_s1_wait_counter_eq_0,
                                       clk,
                                       col_s1_readdata_from_sa,
                                       cpu_0_data_master_address,
                                       cpu_0_data_master_byteenable,
                                       cpu_0_data_master_byteenable_cfi_flash_0_s1,
                                       cpu_0_data_master_byteenable_sdram_0_s1,
                                       cpu_0_data_master_granted_button_pio_s1,
                                       cpu_0_data_master_granted_cfi_flash_0_s1,
                                       cpu_0_data_master_granted_col_s1,
                                       cpu_0_data_master_granted_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_granted_led_pio_s1,
                                       cpu_0_data_master_granted_row_s1,
                                       cpu_0_data_master_granted_sdram_0_s1,
                                       cpu_0_data_master_granted_tft_lcd_data_s1,
                                       cpu_0_data_master_granted_tft_lcd_nrd_s1,
                                       cpu_0_data_master_granted_tft_lcd_nrst_s1,
                                       cpu_0_data_master_granted_tft_lcd_nwr_s1,
                                       cpu_0_data_master_granted_tft_lcd_rs_s1,
                                       cpu_0_data_master_qualified_request_button_pio_s1,
                                       cpu_0_data_master_qualified_request_cfi_flash_0_s1,
                                       cpu_0_data_master_qualified_request_col_s1,
                                       cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_qualified_request_led_pio_s1,
                                       cpu_0_data_master_qualified_request_row_s1,
                                       cpu_0_data_master_qualified_request_sdram_0_s1,
                                       cpu_0_data_master_qualified_request_tft_lcd_data_s1,
                                       cpu_0_data_master_qualified_request_tft_lcd_nrd_s1,
                                       cpu_0_data_master_qualified_request_tft_lcd_nrst_s1,
                                       cpu_0_data_master_qualified_request_tft_lcd_nwr_s1,
                                       cpu_0_data_master_qualified_request_tft_lcd_rs_s1,
                                       cpu_0_data_master_read,
                                       cpu_0_data_master_read_data_valid_button_pio_s1,
                                       cpu_0_data_master_read_data_valid_cfi_flash_0_s1,
                                       cpu_0_data_master_read_data_valid_col_s1,
                                       cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_read_data_valid_led_pio_s1,
                                       cpu_0_data_master_read_data_valid_row_s1,
                                       cpu_0_data_master_read_data_valid_sdram_0_s1,
                                       cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                       cpu_0_data_master_read_data_valid_tft_lcd_data_s1,
                                       cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1,
                                       cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1,
                                       cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1,
                                       cpu_0_data_master_read_data_valid_tft_lcd_rs_s1,
                                       cpu_0_data_master_requests_button_pio_s1,
                                       cpu_0_data_master_requests_cfi_flash_0_s1,
                                       cpu_0_data_master_requests_col_s1,
                                       cpu_0_data_master_requests_cpu_0_jtag_debug_module,
                                       cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave,
                                       cpu_0_data_master_requests_led_pio_s1,
                                       cpu_0_data_master_requests_row_s1,
                                       cpu_0_data_master_requests_sdram_0_s1,
                                       cpu_0_data_master_requests_tft_lcd_data_s1,
                                       cpu_0_data_master_requests_tft_lcd_nrd_s1,
                                       cpu_0_data_master_requests_tft_lcd_nrst_s1,
                                       cpu_0_data_master_requests_tft_lcd_nwr_s1,
                                       cpu_0_data_master_requests_tft_lcd_rs_s1,
                                       cpu_0_data_master_write,
                                       cpu_0_data_master_writedata,
                                       cpu_0_jtag_debug_module_readdata_from_sa,
                                       d1_button_pio_s1_end_xfer,
                                       d1_col_s1_end_xfer,
                                       d1_cpu_0_jtag_debug_module_end_xfer,
                                       d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                       d1_led_pio_s1_end_xfer,
                                       d1_row_s1_end_xfer,
                                       d1_sdram_0_s1_end_xfer,
                                       d1_tft_lcd_data_s1_end_xfer,
                                       d1_tft_lcd_nrd_s1_end_xfer,
                                       d1_tft_lcd_nrst_s1_end_xfer,
                                       d1_tft_lcd_nwr_s1_end_xfer,
                                       d1_tft_lcd_rs_s1_end_xfer,
                                       d1_tri_state_bridge_0_avalon_slave_end_xfer,
                                       incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0,
                                       jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                       jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                       jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                       led_pio_s1_readdata_from_sa,
                                       reset_n,
                                       row_s1_readdata_from_sa,
                                       sdram_0_s1_readdata_from_sa,
                                       sdram_0_s1_waitrequest_from_sa,
                                       tft_lcd_data_s1_readdata_from_sa,
                                       tft_lcd_nrd_s1_readdata_from_sa,
                                       tft_lcd_nrst_s1_readdata_from_sa,
                                       tft_lcd_nwr_s1_readdata_from_sa,
                                       tft_lcd_rs_s1_readdata_from_sa,

                                      // outputs:
                                       cpu_0_data_master_address_to_slave,
                                       cpu_0_data_master_dbs_address,
                                       cpu_0_data_master_dbs_write_16,
                                       cpu_0_data_master_irq,
                                       cpu_0_data_master_latency_counter,
                                       cpu_0_data_master_readdata,
                                       cpu_0_data_master_readdatavalid,
                                       cpu_0_data_master_waitrequest
                                    )
;

  output  [ 24: 0] cpu_0_data_master_address_to_slave;
  output  [  1: 0] cpu_0_data_master_dbs_address;
  output  [ 15: 0] cpu_0_data_master_dbs_write_16;
  output  [ 31: 0] cpu_0_data_master_irq;
  output  [  1: 0] cpu_0_data_master_latency_counter;
  output  [ 31: 0] cpu_0_data_master_readdata;
  output           cpu_0_data_master_readdatavalid;
  output           cpu_0_data_master_waitrequest;
  input            button_pio_s1_irq_from_sa;
  input   [  7: 0] button_pio_s1_readdata_from_sa;
  input            cfi_flash_0_s1_wait_counter_eq_0;
  input            clk;
  input   [  3: 0] col_s1_readdata_from_sa;
  input   [ 24: 0] cpu_0_data_master_address;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1;
  input   [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1;
  input            cpu_0_data_master_granted_button_pio_s1;
  input            cpu_0_data_master_granted_cfi_flash_0_s1;
  input            cpu_0_data_master_granted_col_s1;
  input            cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_granted_led_pio_s1;
  input            cpu_0_data_master_granted_row_s1;
  input            cpu_0_data_master_granted_sdram_0_s1;
  input            cpu_0_data_master_granted_tft_lcd_data_s1;
  input            cpu_0_data_master_granted_tft_lcd_nrd_s1;
  input            cpu_0_data_master_granted_tft_lcd_nrst_s1;
  input            cpu_0_data_master_granted_tft_lcd_nwr_s1;
  input            cpu_0_data_master_granted_tft_lcd_rs_s1;
  input            cpu_0_data_master_qualified_request_button_pio_s1;
  input            cpu_0_data_master_qualified_request_cfi_flash_0_s1;
  input            cpu_0_data_master_qualified_request_col_s1;
  input            cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_qualified_request_led_pio_s1;
  input            cpu_0_data_master_qualified_request_row_s1;
  input            cpu_0_data_master_qualified_request_sdram_0_s1;
  input            cpu_0_data_master_qualified_request_tft_lcd_data_s1;
  input            cpu_0_data_master_qualified_request_tft_lcd_nrd_s1;
  input            cpu_0_data_master_qualified_request_tft_lcd_nrst_s1;
  input            cpu_0_data_master_qualified_request_tft_lcd_nwr_s1;
  input            cpu_0_data_master_qualified_request_tft_lcd_rs_s1;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_button_pio_s1;
  input            cpu_0_data_master_read_data_valid_cfi_flash_0_s1;
  input            cpu_0_data_master_read_data_valid_col_s1;
  input            cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_read_data_valid_led_pio_s1;
  input            cpu_0_data_master_read_data_valid_row_s1;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_read_data_valid_tft_lcd_data_s1;
  input            cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1;
  input            cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1;
  input            cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1;
  input            cpu_0_data_master_read_data_valid_tft_lcd_rs_s1;
  input            cpu_0_data_master_requests_button_pio_s1;
  input            cpu_0_data_master_requests_cfi_flash_0_s1;
  input            cpu_0_data_master_requests_col_s1;
  input            cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  input            cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  input            cpu_0_data_master_requests_led_pio_s1;
  input            cpu_0_data_master_requests_row_s1;
  input            cpu_0_data_master_requests_sdram_0_s1;
  input            cpu_0_data_master_requests_tft_lcd_data_s1;
  input            cpu_0_data_master_requests_tft_lcd_nrd_s1;
  input            cpu_0_data_master_requests_tft_lcd_nrst_s1;
  input            cpu_0_data_master_requests_tft_lcd_nwr_s1;
  input            cpu_0_data_master_requests_tft_lcd_rs_s1;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  input            d1_button_pio_s1_end_xfer;
  input            d1_col_s1_end_xfer;
  input            d1_cpu_0_jtag_debug_module_end_xfer;
  input            d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  input            d1_led_pio_s1_end_xfer;
  input            d1_row_s1_end_xfer;
  input            d1_sdram_0_s1_end_xfer;
  input            d1_tft_lcd_data_s1_end_xfer;
  input            d1_tft_lcd_nrd_s1_end_xfer;
  input            d1_tft_lcd_nrst_s1_end_xfer;
  input            d1_tft_lcd_nwr_s1_end_xfer;
  input            d1_tft_lcd_rs_s1_end_xfer;
  input            d1_tri_state_bridge_0_avalon_slave_end_xfer;
  input   [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0;
  input            jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  input   [  7: 0] led_pio_s1_readdata_from_sa;
  input            reset_n;
  input   [ 15: 0] row_s1_readdata_from_sa;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;
  input   [  7: 0] tft_lcd_data_s1_readdata_from_sa;
  input            tft_lcd_nrd_s1_readdata_from_sa;
  input            tft_lcd_nrst_s1_readdata_from_sa;
  input            tft_lcd_nwr_s1_readdata_from_sa;
  input            tft_lcd_rs_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_0_data_master_address_last_time;
  wire    [ 24: 0] cpu_0_data_master_address_to_slave;
  reg     [  3: 0] cpu_0_data_master_byteenable_last_time;
  reg     [  1: 0] cpu_0_data_master_dbs_address;
  wire    [  1: 0] cpu_0_data_master_dbs_increment;
  reg     [  1: 0] cpu_0_data_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_0_data_master_dbs_rdv_counter_inc;
  wire    [ 15: 0] cpu_0_data_master_dbs_write_16;
  wire    [ 31: 0] cpu_0_data_master_irq;
  wire             cpu_0_data_master_is_granted_some_slave;
  reg     [  1: 0] cpu_0_data_master_latency_counter;
  wire    [  1: 0] cpu_0_data_master_next_dbs_rdv_counter;
  reg              cpu_0_data_master_read_but_no_slave_selected;
  reg              cpu_0_data_master_read_last_time;
  wire    [ 31: 0] cpu_0_data_master_readdata;
  wire             cpu_0_data_master_readdatavalid;
  wire             cpu_0_data_master_run;
  wire             cpu_0_data_master_waitrequest;
  reg              cpu_0_data_master_write_last_time;
  reg     [ 31: 0] cpu_0_data_master_writedata_last_time;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [  1: 0] p1_cpu_0_data_master_latency_counter;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_0_data_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_0_data_master_qualified_request_button_pio_s1 | ~cpu_0_data_master_requests_button_pio_s1) & ((~cpu_0_data_master_qualified_request_button_pio_s1 | ~cpu_0_data_master_read | (1 & ~d1_button_pio_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_button_pio_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_col_s1 | ~cpu_0_data_master_requests_col_s1) & ((~cpu_0_data_master_qualified_request_col_s1 | ~cpu_0_data_master_read | (1 & ~d1_col_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_col_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_requests_cpu_0_jtag_debug_module) & (cpu_0_data_master_granted_cpu_0_jtag_debug_module | ~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module) & ((~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_read | (1 & ~d1_cpu_0_jtag_debug_module_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave) & ((~cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (cpu_0_data_master_read | cpu_0_data_master_write)))) & ((~cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave | ~(cpu_0_data_master_read | cpu_0_data_master_write) | (1 & ~jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa & (cpu_0_data_master_read | cpu_0_data_master_write)))) & 1 & (cpu_0_data_master_qualified_request_led_pio_s1 | ~cpu_0_data_master_requests_led_pio_s1) & ((~cpu_0_data_master_qualified_request_led_pio_s1 | ~cpu_0_data_master_read | (1 & ~d1_led_pio_s1_end_xfer & cpu_0_data_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_0_data_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = ((~cpu_0_data_master_qualified_request_led_pio_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_row_s1 | ~cpu_0_data_master_requests_row_s1) & ((~cpu_0_data_master_qualified_request_row_s1 | ~cpu_0_data_master_read | (1 & ~d1_row_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_row_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_sdram_0_s1 | (cpu_0_data_master_write & !cpu_0_data_master_byteenable_sdram_0_s1 & cpu_0_data_master_dbs_address[1]) | ~cpu_0_data_master_requests_sdram_0_s1) & (cpu_0_data_master_granted_sdram_0_s1 | ~cpu_0_data_master_qualified_request_sdram_0_s1) & ((~cpu_0_data_master_qualified_request_sdram_0_s1 | ~cpu_0_data_master_read | (1 & ~sdram_0_s1_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_sdram_0_s1 | ~cpu_0_data_master_write | (1 & ~sdram_0_s1_waitrequest_from_sa & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_tft_lcd_data_s1 | ~cpu_0_data_master_requests_tft_lcd_data_s1) & (cpu_0_data_master_granted_tft_lcd_data_s1 | ~cpu_0_data_master_qualified_request_tft_lcd_data_s1) & ((~cpu_0_data_master_qualified_request_tft_lcd_data_s1 | ~cpu_0_data_master_read | (1 & ~d1_tft_lcd_data_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_tft_lcd_data_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 | ~cpu_0_data_master_requests_tft_lcd_nrd_s1) & (cpu_0_data_master_granted_tft_lcd_nrd_s1 | ~cpu_0_data_master_qualified_request_tft_lcd_nrd_s1) & ((~cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 | ~cpu_0_data_master_read | (1 & ~d1_tft_lcd_nrd_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 | ~cpu_0_data_master_requests_tft_lcd_nrst_s1) & (cpu_0_data_master_granted_tft_lcd_nrst_s1 | ~cpu_0_data_master_qualified_request_tft_lcd_nrst_s1) & ((~cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 | ~cpu_0_data_master_read | (1 & ~d1_tft_lcd_nrst_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 | ~cpu_0_data_master_requests_tft_lcd_nwr_s1) & (cpu_0_data_master_granted_tft_lcd_nwr_s1 | ~cpu_0_data_master_qualified_request_tft_lcd_nwr_s1) & ((~cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 | ~cpu_0_data_master_read | (1 & ~d1_tft_lcd_nwr_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_tft_lcd_rs_s1 | ~cpu_0_data_master_requests_tft_lcd_rs_s1) & (cpu_0_data_master_granted_tft_lcd_rs_s1 | ~cpu_0_data_master_qualified_request_tft_lcd_rs_s1) & ((~cpu_0_data_master_qualified_request_tft_lcd_rs_s1 | ~cpu_0_data_master_read | (1 & ~d1_tft_lcd_rs_s1_end_xfer & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_tft_lcd_rs_s1 | ~cpu_0_data_master_write | (1 & cpu_0_data_master_write))) & 1 & (cpu_0_data_master_qualified_request_cfi_flash_0_s1 | (cpu_0_data_master_write & !cpu_0_data_master_byteenable_cfi_flash_0_s1 & cpu_0_data_master_dbs_address[1]) | ~cpu_0_data_master_requests_cfi_flash_0_s1) & (cpu_0_data_master_granted_cfi_flash_0_s1 | ~cpu_0_data_master_qualified_request_cfi_flash_0_s1) & ((~cpu_0_data_master_qualified_request_cfi_flash_0_s1 | ~cpu_0_data_master_read | (1 & ((cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer)) & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_read))) & ((~cpu_0_data_master_qualified_request_cfi_flash_0_s1 | ~cpu_0_data_master_write | (1 & ((cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer)) & (cpu_0_data_master_dbs_address[1]) & cpu_0_data_master_write)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_0_data_master_address_to_slave = cpu_0_data_master_address[24 : 0];

  //cpu_0_data_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_but_no_slave_selected <= 0;
      else 
        cpu_0_data_master_read_but_no_slave_selected <= cpu_0_data_master_read & cpu_0_data_master_run & ~cpu_0_data_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_0_data_master_is_granted_some_slave = cpu_0_data_master_granted_button_pio_s1 |
    cpu_0_data_master_granted_col_s1 |
    cpu_0_data_master_granted_cpu_0_jtag_debug_module |
    cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave |
    cpu_0_data_master_granted_led_pio_s1 |
    cpu_0_data_master_granted_row_s1 |
    cpu_0_data_master_granted_sdram_0_s1 |
    cpu_0_data_master_granted_tft_lcd_data_s1 |
    cpu_0_data_master_granted_tft_lcd_nrd_s1 |
    cpu_0_data_master_granted_tft_lcd_nrst_s1 |
    cpu_0_data_master_granted_tft_lcd_nwr_s1 |
    cpu_0_data_master_granted_tft_lcd_rs_s1 |
    cpu_0_data_master_granted_cfi_flash_0_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_0_data_master_readdatavalid = (cpu_0_data_master_read_data_valid_sdram_0_s1 & dbs_rdv_counter_overflow) |
    (cpu_0_data_master_read_data_valid_cfi_flash_0_s1 & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_0_data_master_readdatavalid = cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_button_pio_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_col_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_led_pio_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_row_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_tft_lcd_data_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid |
    cpu_0_data_master_read_data_valid_tft_lcd_rs_s1 |
    cpu_0_data_master_read_but_no_slave_selected |
    pre_flush_cpu_0_data_master_readdatavalid;

  //cpu_0/data_master readdata mux, which is an e_mux
  assign cpu_0_data_master_readdata = ({32 {~(cpu_0_data_master_qualified_request_button_pio_s1 & cpu_0_data_master_read)}} | button_pio_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_col_s1 & cpu_0_data_master_read)}} | col_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module & cpu_0_data_master_read)}} | cpu_0_jtag_debug_module_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read)}} | jtag_uart_0_avalon_jtag_slave_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_led_pio_s1 & cpu_0_data_master_read)}} | led_pio_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_row_s1 & cpu_0_data_master_read)}} | row_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_sdram_0_s1}} | {sdram_0_s1_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_0_data_master_qualified_request_tft_lcd_data_s1 & cpu_0_data_master_read)}} | tft_lcd_data_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 & cpu_0_data_master_read)}} | tft_lcd_nrd_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 & cpu_0_data_master_read)}} | tft_lcd_nrst_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 & cpu_0_data_master_read)}} | tft_lcd_nwr_s1_readdata_from_sa) &
    ({32 {~(cpu_0_data_master_qualified_request_tft_lcd_rs_s1 & cpu_0_data_master_read)}} | tft_lcd_rs_s1_readdata_from_sa) &
    ({32 {~cpu_0_data_master_read_data_valid_cfi_flash_0_s1}} | {incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_0_data_master_waitrequest = ~cpu_0_data_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_latency_counter <= 0;
      else 
        cpu_0_data_master_latency_counter <= p1_cpu_0_data_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_0_data_master_latency_counter = ((cpu_0_data_master_run & cpu_0_data_master_read))? latency_load_value :
    (cpu_0_data_master_latency_counter)? cpu_0_data_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {2 {cpu_0_data_master_requests_cfi_flash_0_s1}} & 2;

  //irq assign, which is an e_assign
  assign cpu_0_data_master_irq = {1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    1'b0,
    button_pio_s1_irq_from_sa,
    jtag_uart_0_avalon_jtag_slave_irq_from_sa};

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (((~0) & cpu_0_data_master_requests_sdram_0_s1 & cpu_0_data_master_write & !cpu_0_data_master_byteenable_sdram_0_s1)) |
    (cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_read & 1 & 1 & ~sdram_0_s1_waitrequest_from_sa) |
    (cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_write & 1 & 1 & ~sdram_0_s1_waitrequest_from_sa) |
    (((~0) & cpu_0_data_master_requests_cfi_flash_0_s1 & cpu_0_data_master_write & !cpu_0_data_master_byteenable_cfi_flash_0_s1)) |
    ((cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_read & 1 & 1 & ({cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer}))) |
    ((cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_write & 1 & 1 & ({cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer})));

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = (cpu_0_data_master_read_data_valid_sdram_0_s1)? sdram_0_s1_readdata_from_sa :
    incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_0_data_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //mux write dbs 1, which is an e_mux
  assign cpu_0_data_master_dbs_write_16 = (cpu_0_data_master_dbs_address[1])? cpu_0_data_master_writedata[31 : 16] :
    (~(cpu_0_data_master_dbs_address[1]))? cpu_0_data_master_writedata[15 : 0] :
    (cpu_0_data_master_dbs_address[1])? cpu_0_data_master_writedata[31 : 16] :
    cpu_0_data_master_writedata[15 : 0];

  //dbs count increment, which is an e_mux
  assign cpu_0_data_master_dbs_increment = (cpu_0_data_master_requests_sdram_0_s1)? 2 :
    (cpu_0_data_master_requests_cfi_flash_0_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_0_data_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_0_data_master_dbs_address + cpu_0_data_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_0_data_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_0_data_master_next_dbs_rdv_counter = cpu_0_data_master_dbs_rdv_counter + cpu_0_data_master_dbs_rdv_counter_inc;

  //cpu_0_data_master_rdv_inc_mux, which is an e_mux
  assign cpu_0_data_master_dbs_rdv_counter_inc = (cpu_0_data_master_read_data_valid_sdram_0_s1)? 2 :
    2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_0_data_master_read_data_valid_sdram_0_s1 |
    cpu_0_data_master_read_data_valid_cfi_flash_0_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_0_data_master_dbs_rdv_counter <= cpu_0_data_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_0_data_master_dbs_rdv_counter[1] & ~cpu_0_data_master_next_dbs_rdv_counter[1];


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0_data_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_address_last_time <= 0;
      else 
        cpu_0_data_master_address_last_time <= cpu_0_data_master_address;
    end


  //cpu_0/data_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_0_data_master_waitrequest & (cpu_0_data_master_read | cpu_0_data_master_write);
    end


  //cpu_0_data_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_address != cpu_0_data_master_address_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_byteenable check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_byteenable_last_time <= 0;
      else 
        cpu_0_data_master_byteenable_last_time <= cpu_0_data_master_byteenable;
    end


  //cpu_0_data_master_byteenable matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_byteenable != cpu_0_data_master_byteenable_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_byteenable did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_last_time <= 0;
      else 
        cpu_0_data_master_read_last_time <= cpu_0_data_master_read;
    end


  //cpu_0_data_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_read != cpu_0_data_master_read_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_read did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_write check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_write_last_time <= 0;
      else 
        cpu_0_data_master_write_last_time <= cpu_0_data_master_write;
    end


  //cpu_0_data_master_write matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_write != cpu_0_data_master_write_last_time))
        begin
          $write("%0d ns: cpu_0_data_master_write did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_data_master_writedata check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_writedata_last_time <= 0;
      else 
        cpu_0_data_master_writedata_last_time <= cpu_0_data_master_writedata;
    end


  //cpu_0_data_master_writedata matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_data_master_writedata != cpu_0_data_master_writedata_last_time) & cpu_0_data_master_write)
        begin
          $write("%0d ns: cpu_0_data_master_writedata did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cpu_0_instruction_master_arbitrator (
                                             // inputs:
                                              cfi_flash_0_s1_wait_counter_eq_0,
                                              clk,
                                              cpu_0_instruction_master_address,
                                              cpu_0_instruction_master_granted_cfi_flash_0_s1,
                                              cpu_0_instruction_master_granted_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_granted_sdram_0_s1,
                                              cpu_0_instruction_master_granted_tft_lcd_data_s1,
                                              cpu_0_instruction_master_granted_tft_lcd_nrd_s1,
                                              cpu_0_instruction_master_granted_tft_lcd_nrst_s1,
                                              cpu_0_instruction_master_granted_tft_lcd_nwr_s1,
                                              cpu_0_instruction_master_granted_tft_lcd_rs_s1,
                                              cpu_0_instruction_master_qualified_request_cfi_flash_0_s1,
                                              cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_qualified_request_sdram_0_s1,
                                              cpu_0_instruction_master_qualified_request_tft_lcd_data_s1,
                                              cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1,
                                              cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1,
                                              cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1,
                                              cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1,
                                              cpu_0_instruction_master_read,
                                              cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1,
                                              cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_read_data_valid_sdram_0_s1,
                                              cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                              cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1,
                                              cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1,
                                              cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1,
                                              cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1,
                                              cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1,
                                              cpu_0_instruction_master_requests_cfi_flash_0_s1,
                                              cpu_0_instruction_master_requests_cpu_0_jtag_debug_module,
                                              cpu_0_instruction_master_requests_sdram_0_s1,
                                              cpu_0_instruction_master_requests_tft_lcd_data_s1,
                                              cpu_0_instruction_master_requests_tft_lcd_nrd_s1,
                                              cpu_0_instruction_master_requests_tft_lcd_nrst_s1,
                                              cpu_0_instruction_master_requests_tft_lcd_nwr_s1,
                                              cpu_0_instruction_master_requests_tft_lcd_rs_s1,
                                              cpu_0_jtag_debug_module_readdata_from_sa,
                                              d1_cpu_0_jtag_debug_module_end_xfer,
                                              d1_sdram_0_s1_end_xfer,
                                              d1_tft_lcd_data_s1_end_xfer,
                                              d1_tft_lcd_nrd_s1_end_xfer,
                                              d1_tft_lcd_nrst_s1_end_xfer,
                                              d1_tft_lcd_nwr_s1_end_xfer,
                                              d1_tft_lcd_rs_s1_end_xfer,
                                              d1_tri_state_bridge_0_avalon_slave_end_xfer,
                                              incoming_data_to_and_from_the_cfi_flash_0,
                                              reset_n,
                                              sdram_0_s1_readdata_from_sa,
                                              sdram_0_s1_waitrequest_from_sa,
                                              tft_lcd_data_s1_readdata_from_sa,
                                              tft_lcd_nrd_s1_readdata_from_sa,
                                              tft_lcd_nrst_s1_readdata_from_sa,
                                              tft_lcd_nwr_s1_readdata_from_sa,
                                              tft_lcd_rs_s1_readdata_from_sa,

                                             // outputs:
                                              cpu_0_instruction_master_address_to_slave,
                                              cpu_0_instruction_master_dbs_address,
                                              cpu_0_instruction_master_latency_counter,
                                              cpu_0_instruction_master_readdata,
                                              cpu_0_instruction_master_readdatavalid,
                                              cpu_0_instruction_master_waitrequest
                                           )
;

  output  [ 24: 0] cpu_0_instruction_master_address_to_slave;
  output  [  1: 0] cpu_0_instruction_master_dbs_address;
  output  [  1: 0] cpu_0_instruction_master_latency_counter;
  output  [ 31: 0] cpu_0_instruction_master_readdata;
  output           cpu_0_instruction_master_readdatavalid;
  output           cpu_0_instruction_master_waitrequest;
  input            cfi_flash_0_s1_wait_counter_eq_0;
  input            clk;
  input   [ 24: 0] cpu_0_instruction_master_address;
  input            cpu_0_instruction_master_granted_cfi_flash_0_s1;
  input            cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_granted_sdram_0_s1;
  input            cpu_0_instruction_master_granted_tft_lcd_data_s1;
  input            cpu_0_instruction_master_granted_tft_lcd_nrd_s1;
  input            cpu_0_instruction_master_granted_tft_lcd_nrst_s1;
  input            cpu_0_instruction_master_granted_tft_lcd_nwr_s1;
  input            cpu_0_instruction_master_granted_tft_lcd_rs_s1;
  input            cpu_0_instruction_master_qualified_request_cfi_flash_0_s1;
  input            cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_qualified_request_sdram_0_s1;
  input            cpu_0_instruction_master_qualified_request_tft_lcd_data_s1;
  input            cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1;
  input            cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1;
  input            cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1;
  input            cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1;
  input            cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1;
  input            cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1;
  input            cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1;
  input            cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1;
  input            cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1;
  input            cpu_0_instruction_master_requests_cfi_flash_0_s1;
  input            cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  input            cpu_0_instruction_master_requests_sdram_0_s1;
  input            cpu_0_instruction_master_requests_tft_lcd_data_s1;
  input            cpu_0_instruction_master_requests_tft_lcd_nrd_s1;
  input            cpu_0_instruction_master_requests_tft_lcd_nrst_s1;
  input            cpu_0_instruction_master_requests_tft_lcd_nwr_s1;
  input            cpu_0_instruction_master_requests_tft_lcd_rs_s1;
  input   [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  input            d1_cpu_0_jtag_debug_module_end_xfer;
  input            d1_sdram_0_s1_end_xfer;
  input            d1_tft_lcd_data_s1_end_xfer;
  input            d1_tft_lcd_nrd_s1_end_xfer;
  input            d1_tft_lcd_nrst_s1_end_xfer;
  input            d1_tft_lcd_nwr_s1_end_xfer;
  input            d1_tft_lcd_rs_s1_end_xfer;
  input            d1_tri_state_bridge_0_avalon_slave_end_xfer;
  input   [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata_from_sa;
  input            sdram_0_s1_waitrequest_from_sa;
  input   [  7: 0] tft_lcd_data_s1_readdata_from_sa;
  input            tft_lcd_nrd_s1_readdata_from_sa;
  input            tft_lcd_nrst_s1_readdata_from_sa;
  input            tft_lcd_nwr_s1_readdata_from_sa;
  input            tft_lcd_rs_s1_readdata_from_sa;

  reg              active_and_waiting_last_time;
  reg     [ 24: 0] cpu_0_instruction_master_address_last_time;
  wire    [ 24: 0] cpu_0_instruction_master_address_to_slave;
  reg     [  1: 0] cpu_0_instruction_master_dbs_address;
  wire    [  1: 0] cpu_0_instruction_master_dbs_increment;
  reg     [  1: 0] cpu_0_instruction_master_dbs_rdv_counter;
  wire    [  1: 0] cpu_0_instruction_master_dbs_rdv_counter_inc;
  wire             cpu_0_instruction_master_is_granted_some_slave;
  reg     [  1: 0] cpu_0_instruction_master_latency_counter;
  wire    [  1: 0] cpu_0_instruction_master_next_dbs_rdv_counter;
  reg              cpu_0_instruction_master_read_but_no_slave_selected;
  reg              cpu_0_instruction_master_read_last_time;
  wire    [ 31: 0] cpu_0_instruction_master_readdata;
  wire             cpu_0_instruction_master_readdatavalid;
  wire             cpu_0_instruction_master_run;
  wire             cpu_0_instruction_master_waitrequest;
  wire             dbs_count_enable;
  wire             dbs_counter_overflow;
  reg     [ 15: 0] dbs_latent_16_reg_segment_0;
  wire             dbs_rdv_count_enable;
  wire             dbs_rdv_counter_overflow;
  wire    [  1: 0] latency_load_value;
  wire    [  1: 0] next_dbs_address;
  wire    [  1: 0] p1_cpu_0_instruction_master_latency_counter;
  wire    [ 15: 0] p1_dbs_latent_16_reg_segment_0;
  wire             pre_dbs_count_enable;
  wire             pre_flush_cpu_0_instruction_master_readdatavalid;
  wire             r_0;
  wire             r_1;
  wire             r_2;
  //r_0 master_run cascaded wait assignment, which is an e_assign
  assign r_0 = 1 & (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_requests_cpu_0_jtag_debug_module) & (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module) & ((~cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module | ~cpu_0_instruction_master_read | (1 & ~d1_cpu_0_jtag_debug_module_end_xfer & cpu_0_instruction_master_read)));

  //cascaded wait assignment, which is an e_assign
  assign cpu_0_instruction_master_run = r_0 & r_1 & r_2;

  //r_1 master_run cascaded wait assignment, which is an e_assign
  assign r_1 = 1 & (cpu_0_instruction_master_qualified_request_sdram_0_s1 | ~cpu_0_instruction_master_requests_sdram_0_s1) & (cpu_0_instruction_master_granted_sdram_0_s1 | ~cpu_0_instruction_master_qualified_request_sdram_0_s1) & ((~cpu_0_instruction_master_qualified_request_sdram_0_s1 | ~cpu_0_instruction_master_read | (1 & ~sdram_0_s1_waitrequest_from_sa & (cpu_0_instruction_master_dbs_address[1]) & cpu_0_instruction_master_read))) & 1 & (cpu_0_instruction_master_qualified_request_tft_lcd_data_s1 | ~cpu_0_instruction_master_requests_tft_lcd_data_s1) & (cpu_0_instruction_master_granted_tft_lcd_data_s1 | ~cpu_0_instruction_master_qualified_request_tft_lcd_data_s1) & ((~cpu_0_instruction_master_qualified_request_tft_lcd_data_s1 | ~cpu_0_instruction_master_read | (1 & ~d1_tft_lcd_data_s1_end_xfer & cpu_0_instruction_master_read))) & 1 & (cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1 | ~cpu_0_instruction_master_requests_tft_lcd_nrd_s1) & (cpu_0_instruction_master_granted_tft_lcd_nrd_s1 | ~cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1) & ((~cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1 | ~cpu_0_instruction_master_read | (1 & ~d1_tft_lcd_nrd_s1_end_xfer & cpu_0_instruction_master_read)));

  //r_2 master_run cascaded wait assignment, which is an e_assign
  assign r_2 = 1 & (cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1 | ~cpu_0_instruction_master_requests_tft_lcd_nrst_s1) & (cpu_0_instruction_master_granted_tft_lcd_nrst_s1 | ~cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1) & ((~cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1 | ~cpu_0_instruction_master_read | (1 & ~d1_tft_lcd_nrst_s1_end_xfer & cpu_0_instruction_master_read))) & 1 & (cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1 | ~cpu_0_instruction_master_requests_tft_lcd_nwr_s1) & (cpu_0_instruction_master_granted_tft_lcd_nwr_s1 | ~cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1) & ((~cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1 | ~cpu_0_instruction_master_read | (1 & ~d1_tft_lcd_nwr_s1_end_xfer & cpu_0_instruction_master_read))) & 1 & (cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1 | ~cpu_0_instruction_master_requests_tft_lcd_rs_s1) & (cpu_0_instruction_master_granted_tft_lcd_rs_s1 | ~cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1) & ((~cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1 | ~cpu_0_instruction_master_read | (1 & ~d1_tft_lcd_rs_s1_end_xfer & cpu_0_instruction_master_read))) & 1 & (cpu_0_instruction_master_qualified_request_cfi_flash_0_s1 | ~cpu_0_instruction_master_requests_cfi_flash_0_s1) & (cpu_0_instruction_master_granted_cfi_flash_0_s1 | ~cpu_0_instruction_master_qualified_request_cfi_flash_0_s1) & ((~cpu_0_instruction_master_qualified_request_cfi_flash_0_s1 | ~cpu_0_instruction_master_read | (1 & ((cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer)) & (cpu_0_instruction_master_dbs_address[1]) & cpu_0_instruction_master_read)));

  //optimize select-logic by passing only those address bits which matter.
  assign cpu_0_instruction_master_address_to_slave = cpu_0_instruction_master_address[24 : 0];

  //cpu_0_instruction_master_read_but_no_slave_selected assignment, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_but_no_slave_selected <= 0;
      else 
        cpu_0_instruction_master_read_but_no_slave_selected <= cpu_0_instruction_master_read & cpu_0_instruction_master_run & ~cpu_0_instruction_master_is_granted_some_slave;
    end


  //some slave is getting selected, which is an e_mux
  assign cpu_0_instruction_master_is_granted_some_slave = cpu_0_instruction_master_granted_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_granted_sdram_0_s1 |
    cpu_0_instruction_master_granted_tft_lcd_data_s1 |
    cpu_0_instruction_master_granted_tft_lcd_nrd_s1 |
    cpu_0_instruction_master_granted_tft_lcd_nrst_s1 |
    cpu_0_instruction_master_granted_tft_lcd_nwr_s1 |
    cpu_0_instruction_master_granted_tft_lcd_rs_s1 |
    cpu_0_instruction_master_granted_cfi_flash_0_s1;

  //latent slave read data valids which may be flushed, which is an e_mux
  assign pre_flush_cpu_0_instruction_master_readdatavalid = (cpu_0_instruction_master_read_data_valid_sdram_0_s1 & dbs_rdv_counter_overflow) |
    (cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1 & dbs_rdv_counter_overflow);

  //latent slave read data valid which is not flushed, which is an e_mux
  assign cpu_0_instruction_master_readdatavalid = cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1 |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1 |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1 |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1 |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid |
    cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1 |
    cpu_0_instruction_master_read_but_no_slave_selected |
    pre_flush_cpu_0_instruction_master_readdatavalid;

  //cpu_0/instruction_master readdata mux, which is an e_mux
  assign cpu_0_instruction_master_readdata = ({32 {~(cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module & cpu_0_instruction_master_read)}} | cpu_0_jtag_debug_module_readdata_from_sa) &
    ({32 {~cpu_0_instruction_master_read_data_valid_sdram_0_s1}} | {sdram_0_s1_readdata_from_sa[15 : 0],
    dbs_latent_16_reg_segment_0}) &
    ({32 {~(cpu_0_instruction_master_qualified_request_tft_lcd_data_s1 & cpu_0_instruction_master_read)}} | tft_lcd_data_s1_readdata_from_sa) &
    ({32 {~(cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1 & cpu_0_instruction_master_read)}} | tft_lcd_nrd_s1_readdata_from_sa) &
    ({32 {~(cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1 & cpu_0_instruction_master_read)}} | tft_lcd_nrst_s1_readdata_from_sa) &
    ({32 {~(cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1 & cpu_0_instruction_master_read)}} | tft_lcd_nwr_s1_readdata_from_sa) &
    ({32 {~(cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1 & cpu_0_instruction_master_read)}} | tft_lcd_rs_s1_readdata_from_sa) &
    ({32 {~cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1}} | {incoming_data_to_and_from_the_cfi_flash_0[15 : 0],
    dbs_latent_16_reg_segment_0});

  //actual waitrequest port, which is an e_assign
  assign cpu_0_instruction_master_waitrequest = ~cpu_0_instruction_master_run;

  //latent max counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_latency_counter <= 0;
      else 
        cpu_0_instruction_master_latency_counter <= p1_cpu_0_instruction_master_latency_counter;
    end


  //latency counter load mux, which is an e_mux
  assign p1_cpu_0_instruction_master_latency_counter = ((cpu_0_instruction_master_run & cpu_0_instruction_master_read))? latency_load_value :
    (cpu_0_instruction_master_latency_counter)? cpu_0_instruction_master_latency_counter - 1 :
    0;

  //read latency load values, which is an e_mux
  assign latency_load_value = {2 {cpu_0_instruction_master_requests_cfi_flash_0_s1}} & 2;

  //input to latent dbs-16 stored 0, which is an e_mux
  assign p1_dbs_latent_16_reg_segment_0 = (cpu_0_instruction_master_read_data_valid_sdram_0_s1)? sdram_0_s1_readdata_from_sa :
    incoming_data_to_and_from_the_cfi_flash_0;

  //dbs register for latent dbs-16 segment 0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          dbs_latent_16_reg_segment_0 <= 0;
      else if (dbs_rdv_count_enable & ((cpu_0_instruction_master_dbs_rdv_counter[1]) == 0))
          dbs_latent_16_reg_segment_0 <= p1_dbs_latent_16_reg_segment_0;
    end


  //dbs count increment, which is an e_mux
  assign cpu_0_instruction_master_dbs_increment = (cpu_0_instruction_master_requests_sdram_0_s1)? 2 :
    (cpu_0_instruction_master_requests_cfi_flash_0_s1)? 2 :
    0;

  //dbs counter overflow, which is an e_assign
  assign dbs_counter_overflow = cpu_0_instruction_master_dbs_address[1] & !(next_dbs_address[1]);

  //next master address, which is an e_assign
  assign next_dbs_address = cpu_0_instruction_master_dbs_address + cpu_0_instruction_master_dbs_increment;

  //dbs count enable, which is an e_mux
  assign dbs_count_enable = pre_dbs_count_enable;

  //dbs counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_dbs_address <= 0;
      else if (dbs_count_enable)
          cpu_0_instruction_master_dbs_address <= next_dbs_address;
    end


  //p1 dbs rdv counter, which is an e_assign
  assign cpu_0_instruction_master_next_dbs_rdv_counter = cpu_0_instruction_master_dbs_rdv_counter + cpu_0_instruction_master_dbs_rdv_counter_inc;

  //cpu_0_instruction_master_rdv_inc_mux, which is an e_mux
  assign cpu_0_instruction_master_dbs_rdv_counter_inc = (cpu_0_instruction_master_read_data_valid_sdram_0_s1)? 2 :
    2;

  //master any slave rdv, which is an e_mux
  assign dbs_rdv_count_enable = cpu_0_instruction_master_read_data_valid_sdram_0_s1 |
    cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1;

  //dbs rdv counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_dbs_rdv_counter <= 0;
      else if (dbs_rdv_count_enable)
          cpu_0_instruction_master_dbs_rdv_counter <= cpu_0_instruction_master_next_dbs_rdv_counter;
    end


  //dbs rdv counter overflow, which is an e_assign
  assign dbs_rdv_counter_overflow = cpu_0_instruction_master_dbs_rdv_counter[1] & ~cpu_0_instruction_master_next_dbs_rdv_counter[1];

  //pre dbs count enable, which is an e_mux
  assign pre_dbs_count_enable = (cpu_0_instruction_master_granted_sdram_0_s1 & cpu_0_instruction_master_read & 1 & 1 & ~sdram_0_s1_waitrequest_from_sa) |
    ((cpu_0_instruction_master_granted_cfi_flash_0_s1 & cpu_0_instruction_master_read & 1 & 1 & ({cfi_flash_0_s1_wait_counter_eq_0 & ~d1_tri_state_bridge_0_avalon_slave_end_xfer})));


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //cpu_0_instruction_master_address check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_address_last_time <= 0;
      else 
        cpu_0_instruction_master_address_last_time <= cpu_0_instruction_master_address;
    end


  //cpu_0/instruction_master waited last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          active_and_waiting_last_time <= 0;
      else 
        active_and_waiting_last_time <= cpu_0_instruction_master_waitrequest & (cpu_0_instruction_master_read);
    end


  //cpu_0_instruction_master_address matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_instruction_master_address != cpu_0_instruction_master_address_last_time))
        begin
          $write("%0d ns: cpu_0_instruction_master_address did not heed wait!!!", $time);
          $stop;
        end
    end


  //cpu_0_instruction_master_read check against wait, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_last_time <= 0;
      else 
        cpu_0_instruction_master_read_last_time <= cpu_0_instruction_master_read;
    end


  //cpu_0_instruction_master_read matches last port_name, which is an e_process
  always @(posedge clk)
    begin
      if (active_and_waiting_last_time & (cpu_0_instruction_master_read != cpu_0_instruction_master_read_last_time))
        begin
          $write("%0d ns: cpu_0_instruction_master_read did not heed wait!!!", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module jtag_uart_0_avalon_jtag_slave_arbitrator (
                                                  // inputs:
                                                   clk,
                                                   cpu_0_data_master_address_to_slave,
                                                   cpu_0_data_master_latency_counter,
                                                   cpu_0_data_master_read,
                                                   cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                                   cpu_0_data_master_write,
                                                   cpu_0_data_master_writedata,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable,
                                                   jtag_uart_0_avalon_jtag_slave_irq,
                                                   jtag_uart_0_avalon_jtag_slave_readdata,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest,
                                                   reset_n,

                                                  // outputs:
                                                   cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave,
                                                   cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave,
                                                   d1_jtag_uart_0_avalon_jtag_slave_end_xfer,
                                                   jtag_uart_0_avalon_jtag_slave_address,
                                                   jtag_uart_0_avalon_jtag_slave_chipselect,
                                                   jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_irq_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_read_n,
                                                   jtag_uart_0_avalon_jtag_slave_readdata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_reset_n,
                                                   jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa,
                                                   jtag_uart_0_avalon_jtag_slave_write_n,
                                                   jtag_uart_0_avalon_jtag_slave_writedata
                                                )
;

  output           cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  output           cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  output           d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  output           jtag_uart_0_avalon_jtag_slave_address;
  output           jtag_uart_0_avalon_jtag_slave_chipselect;
  output           jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_read_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_reset_n;
  output           jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  output           jtag_uart_0_avalon_jtag_slave_write_n;
  output  [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input            jtag_uart_0_avalon_jtag_slave_dataavailable;
  input            jtag_uart_0_avalon_jtag_slave_irq;
  input   [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  input            jtag_uart_0_avalon_jtag_slave_readyfordata;
  input            jtag_uart_0_avalon_jtag_slave_waitrequest;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_saved_grant_jtag_uart_0_avalon_jtag_slave;
  reg              d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_allgrants;
  wire             jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant;
  wire             jtag_uart_0_avalon_jtag_slave_any_continuerequest;
  wire             jtag_uart_0_avalon_jtag_slave_arb_counter_enable;
  reg     [  1: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter;
  wire    [  1: 0] jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
  wire    [  1: 0] jtag_uart_0_avalon_jtag_slave_arb_share_set_values;
  wire             jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal;
  wire             jtag_uart_0_avalon_jtag_slave_begins_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             jtag_uart_0_avalon_jtag_slave_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_grant_vector;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_master_qreq_vector;
  wire             jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  reg              jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  reg              jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable;
  wire             jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2;
  wire             jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_read;
  wire             jtag_uart_0_avalon_jtag_slave_waits_for_write;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire    [ 24: 0] shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master;
  wire             wait_for_jtag_uart_0_avalon_jtag_slave_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  assign jtag_uart_0_avalon_jtag_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave));
  //assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readdata_from_sa = jtag_uart_0_avalon_jtag_slave_readdata;

  assign cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave = ({cpu_0_data_master_address_to_slave[24 : 3] , 3'b0} == 25'h18010e0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa = jtag_uart_0_avalon_jtag_slave_dataavailable;

  //assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa = jtag_uart_0_avalon_jtag_slave_readyfordata;

  //assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa = jtag_uart_0_avalon_jtag_slave_waitrequest;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter set values, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_arb_share_set_values = 1;

  //jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;

  //jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant = 0;

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value = jtag_uart_0_avalon_jtag_slave_firsttransfer ? (jtag_uart_0_avalon_jtag_slave_arb_share_set_values - 1) : |jtag_uart_0_avalon_jtag_slave_arb_share_counter ? (jtag_uart_0_avalon_jtag_slave_arb_share_counter - 1) : 0;

  //jtag_uart_0_avalon_jtag_slave_allgrants all slave grants, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_allgrants = |jtag_uart_0_avalon_jtag_slave_grant_vector;

  //jtag_uart_0_avalon_jtag_slave_end_xfer assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_end_xfer = ~(jtag_uart_0_avalon_jtag_slave_waits_for_read | jtag_uart_0_avalon_jtag_slave_waits_for_write);

  //end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave = jtag_uart_0_avalon_jtag_slave_end_xfer & (~jtag_uart_0_avalon_jtag_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & jtag_uart_0_avalon_jtag_slave_allgrants) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests);

  //jtag_uart_0_avalon_jtag_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= 0;
      else if (jtag_uart_0_avalon_jtag_slave_arb_counter_enable)
          jtag_uart_0_avalon_jtag_slave_arb_share_counter <= jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= 0;
      else if ((|jtag_uart_0_avalon_jtag_slave_master_qreq_vector & end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave) | (end_xfer_arb_share_counter_term_jtag_uart_0_avalon_jtag_slave & ~jtag_uart_0_avalon_jtag_slave_non_bursting_master_requests))
          jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable <= |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master jtag_uart_0/avalon_jtag_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 = |jtag_uart_0_avalon_jtag_slave_arb_share_counter_next_value;

  //cpu_0/data_master jtag_uart_0/avalon_jtag_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //jtag_uart_0_avalon_jtag_slave_any_continuerequest at least one master continues requesting, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave, which is an e_mux
  assign cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read & ~jtag_uart_0_avalon_jtag_slave_waits_for_read;

  //jtag_uart_0_avalon_jtag_slave_writedata mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;

  //cpu_0/data_master saved-grant jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign cpu_0_data_master_saved_grant_jtag_uart_0_avalon_jtag_slave = cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;

  //allow new arb cycle for jtag_uart_0/avalon_jtag_slave, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign jtag_uart_0_avalon_jtag_slave_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign jtag_uart_0_avalon_jtag_slave_master_qreq_vector = 1;

  //jtag_uart_0_avalon_jtag_slave_reset_n assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_reset_n = reset_n;

  assign jtag_uart_0_avalon_jtag_slave_chipselect = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  //jtag_uart_0_avalon_jtag_slave_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_firsttransfer = jtag_uart_0_avalon_jtag_slave_begins_xfer ? jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer : jtag_uart_0_avalon_jtag_slave_reg_firsttransfer;

  //jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer = ~(jtag_uart_0_avalon_jtag_slave_slavearbiterlockenable & jtag_uart_0_avalon_jtag_slave_any_continuerequest);

  //jtag_uart_0_avalon_jtag_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= 1'b1;
      else if (jtag_uart_0_avalon_jtag_slave_begins_xfer)
          jtag_uart_0_avalon_jtag_slave_reg_firsttransfer <= jtag_uart_0_avalon_jtag_slave_unreg_firsttransfer;
    end


  //jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_beginbursttransfer_internal = jtag_uart_0_avalon_jtag_slave_begins_xfer;

  //~jtag_uart_0_avalon_jtag_slave_read_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_read_n = ~(cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read);

  //~jtag_uart_0_avalon_jtag_slave_write_n assignment, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_write_n = ~(cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_write);

  assign shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //jtag_uart_0_avalon_jtag_slave_address mux, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_address = shifted_address_to_jtag_uart_0_avalon_jtag_slave_from_cpu_0_data_master >> 2;

  //d1_jtag_uart_0_avalon_jtag_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= 1;
      else 
        d1_jtag_uart_0_avalon_jtag_slave_end_xfer <= jtag_uart_0_avalon_jtag_slave_end_xfer;
    end


  //jtag_uart_0_avalon_jtag_slave_waits_for_read in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_read = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_read_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_read_cycle = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = jtag_uart_0_avalon_jtag_slave_in_a_read_cycle;

  //jtag_uart_0_avalon_jtag_slave_waits_for_write in a cycle, which is an e_mux
  assign jtag_uart_0_avalon_jtag_slave_waits_for_write = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle & jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;

  //jtag_uart_0_avalon_jtag_slave_in_a_write_cycle assignment, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_in_a_write_cycle = cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = jtag_uart_0_avalon_jtag_slave_in_a_write_cycle;

  assign wait_for_jtag_uart_0_avalon_jtag_slave_counter = 0;
  //assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign jtag_uart_0_avalon_jtag_slave_irq_from_sa = jtag_uart_0_avalon_jtag_slave_irq;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //jtag_uart_0/avalon_jtag_slave enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module led_pio_s1_arbitrator (
                               // inputs:
                                clk,
                                cpu_0_data_master_address_to_slave,
                                cpu_0_data_master_byteenable,
                                cpu_0_data_master_latency_counter,
                                cpu_0_data_master_read,
                                cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                cpu_0_data_master_write,
                                cpu_0_data_master_writedata,
                                led_pio_s1_readdata,
                                reset_n,

                               // outputs:
                                cpu_0_data_master_granted_led_pio_s1,
                                cpu_0_data_master_qualified_request_led_pio_s1,
                                cpu_0_data_master_read_data_valid_led_pio_s1,
                                cpu_0_data_master_requests_led_pio_s1,
                                d1_led_pio_s1_end_xfer,
                                led_pio_s1_address,
                                led_pio_s1_chipselect,
                                led_pio_s1_readdata_from_sa,
                                led_pio_s1_reset_n,
                                led_pio_s1_write_n,
                                led_pio_s1_writedata
                             )
;

  output           cpu_0_data_master_granted_led_pio_s1;
  output           cpu_0_data_master_qualified_request_led_pio_s1;
  output           cpu_0_data_master_read_data_valid_led_pio_s1;
  output           cpu_0_data_master_requests_led_pio_s1;
  output           d1_led_pio_s1_end_xfer;
  output  [  1: 0] led_pio_s1_address;
  output           led_pio_s1_chipselect;
  output  [  7: 0] led_pio_s1_readdata_from_sa;
  output           led_pio_s1_reset_n;
  output           led_pio_s1_write_n;
  output  [  7: 0] led_pio_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [  7: 0] led_pio_s1_readdata;
  input            reset_n;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_led_pio_s1;
  wire             cpu_0_data_master_qualified_request_led_pio_s1;
  wire             cpu_0_data_master_read_data_valid_led_pio_s1;
  wire             cpu_0_data_master_requests_led_pio_s1;
  wire             cpu_0_data_master_saved_grant_led_pio_s1;
  reg              d1_led_pio_s1_end_xfer;
  reg              d1_reasons_to_wait;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_led_pio_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_allgrants;
  wire             led_pio_s1_allow_new_arb_cycle;
  wire             led_pio_s1_any_bursting_master_saved_grant;
  wire             led_pio_s1_any_continuerequest;
  wire             led_pio_s1_arb_counter_enable;
  reg     [  1: 0] led_pio_s1_arb_share_counter;
  wire    [  1: 0] led_pio_s1_arb_share_counter_next_value;
  wire    [  1: 0] led_pio_s1_arb_share_set_values;
  wire             led_pio_s1_beginbursttransfer_internal;
  wire             led_pio_s1_begins_xfer;
  wire             led_pio_s1_chipselect;
  wire             led_pio_s1_end_xfer;
  wire             led_pio_s1_firsttransfer;
  wire             led_pio_s1_grant_vector;
  wire             led_pio_s1_in_a_read_cycle;
  wire             led_pio_s1_in_a_write_cycle;
  wire             led_pio_s1_master_qreq_vector;
  wire             led_pio_s1_non_bursting_master_requests;
  wire             led_pio_s1_pretend_byte_enable;
  wire    [  7: 0] led_pio_s1_readdata_from_sa;
  reg              led_pio_s1_reg_firsttransfer;
  wire             led_pio_s1_reset_n;
  reg              led_pio_s1_slavearbiterlockenable;
  wire             led_pio_s1_slavearbiterlockenable2;
  wire             led_pio_s1_unreg_firsttransfer;
  wire             led_pio_s1_waits_for_read;
  wire             led_pio_s1_waits_for_write;
  wire             led_pio_s1_write_n;
  wire    [  7: 0] led_pio_s1_writedata;
  wire    [ 24: 0] shifted_address_to_led_pio_s1_from_cpu_0_data_master;
  wire             wait_for_led_pio_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~led_pio_s1_end_xfer;
    end


  assign led_pio_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_led_pio_s1));
  //assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign led_pio_s1_readdata_from_sa = led_pio_s1_readdata;

  assign cpu_0_data_master_requests_led_pio_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801060) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //led_pio_s1_arb_share_counter set values, which is an e_mux
  assign led_pio_s1_arb_share_set_values = 1;

  //led_pio_s1_non_bursting_master_requests mux, which is an e_mux
  assign led_pio_s1_non_bursting_master_requests = cpu_0_data_master_requests_led_pio_s1;

  //led_pio_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign led_pio_s1_any_bursting_master_saved_grant = 0;

  //led_pio_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign led_pio_s1_arb_share_counter_next_value = led_pio_s1_firsttransfer ? (led_pio_s1_arb_share_set_values - 1) : |led_pio_s1_arb_share_counter ? (led_pio_s1_arb_share_counter - 1) : 0;

  //led_pio_s1_allgrants all slave grants, which is an e_mux
  assign led_pio_s1_allgrants = |led_pio_s1_grant_vector;

  //led_pio_s1_end_xfer assignment, which is an e_assign
  assign led_pio_s1_end_xfer = ~(led_pio_s1_waits_for_read | led_pio_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_led_pio_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_led_pio_s1 = led_pio_s1_end_xfer & (~led_pio_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //led_pio_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign led_pio_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_led_pio_s1 & led_pio_s1_allgrants) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests);

  //led_pio_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_arb_share_counter <= 0;
      else if (led_pio_s1_arb_counter_enable)
          led_pio_s1_arb_share_counter <= led_pio_s1_arb_share_counter_next_value;
    end


  //led_pio_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_slavearbiterlockenable <= 0;
      else if ((|led_pio_s1_master_qreq_vector & end_xfer_arb_share_counter_term_led_pio_s1) | (end_xfer_arb_share_counter_term_led_pio_s1 & ~led_pio_s1_non_bursting_master_requests))
          led_pio_s1_slavearbiterlockenable <= |led_pio_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master led_pio/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = led_pio_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //led_pio_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign led_pio_s1_slavearbiterlockenable2 = |led_pio_s1_arb_share_counter_next_value;

  //cpu_0/data_master led_pio/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = led_pio_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //led_pio_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign led_pio_s1_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_led_pio_s1 = cpu_0_data_master_requests_led_pio_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_led_pio_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_led_pio_s1 = cpu_0_data_master_granted_led_pio_s1 & cpu_0_data_master_read & ~led_pio_s1_waits_for_read;

  //led_pio_s1_writedata mux, which is an e_mux
  assign led_pio_s1_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_led_pio_s1 = cpu_0_data_master_qualified_request_led_pio_s1;

  //cpu_0/data_master saved-grant led_pio/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_led_pio_s1 = cpu_0_data_master_requests_led_pio_s1;

  //allow new arb cycle for led_pio/s1, which is an e_assign
  assign led_pio_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign led_pio_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign led_pio_s1_master_qreq_vector = 1;

  //led_pio_s1_reset_n assignment, which is an e_assign
  assign led_pio_s1_reset_n = reset_n;

  assign led_pio_s1_chipselect = cpu_0_data_master_granted_led_pio_s1;
  //led_pio_s1_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_firsttransfer = led_pio_s1_begins_xfer ? led_pio_s1_unreg_firsttransfer : led_pio_s1_reg_firsttransfer;

  //led_pio_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign led_pio_s1_unreg_firsttransfer = ~(led_pio_s1_slavearbiterlockenable & led_pio_s1_any_continuerequest);

  //led_pio_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          led_pio_s1_reg_firsttransfer <= 1'b1;
      else if (led_pio_s1_begins_xfer)
          led_pio_s1_reg_firsttransfer <= led_pio_s1_unreg_firsttransfer;
    end


  //led_pio_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign led_pio_s1_beginbursttransfer_internal = led_pio_s1_begins_xfer;

  //~led_pio_s1_write_n assignment, which is an e_mux
  assign led_pio_s1_write_n = ~(((cpu_0_data_master_granted_led_pio_s1 & cpu_0_data_master_write)) & led_pio_s1_pretend_byte_enable);

  assign shifted_address_to_led_pio_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //led_pio_s1_address mux, which is an e_mux
  assign led_pio_s1_address = shifted_address_to_led_pio_s1_from_cpu_0_data_master >> 2;

  //d1_led_pio_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_led_pio_s1_end_xfer <= 1;
      else 
        d1_led_pio_s1_end_xfer <= led_pio_s1_end_xfer;
    end


  //led_pio_s1_waits_for_read in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_read = led_pio_s1_in_a_read_cycle & led_pio_s1_begins_xfer;

  //led_pio_s1_in_a_read_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_read_cycle = cpu_0_data_master_granted_led_pio_s1 & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = led_pio_s1_in_a_read_cycle;

  //led_pio_s1_waits_for_write in a cycle, which is an e_mux
  assign led_pio_s1_waits_for_write = led_pio_s1_in_a_write_cycle & 0;

  //led_pio_s1_in_a_write_cycle assignment, which is an e_assign
  assign led_pio_s1_in_a_write_cycle = cpu_0_data_master_granted_led_pio_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = led_pio_s1_in_a_write_cycle;

  assign wait_for_led_pio_s1_counter = 0;
  //led_pio_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  assign led_pio_s1_pretend_byte_enable = (cpu_0_data_master_granted_led_pio_s1)? cpu_0_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //led_pio/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module row_s1_arbitrator (
                           // inputs:
                            clk,
                            cpu_0_data_master_address_to_slave,
                            cpu_0_data_master_latency_counter,
                            cpu_0_data_master_read,
                            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                            cpu_0_data_master_write,
                            cpu_0_data_master_writedata,
                            reset_n,
                            row_s1_readdata,

                           // outputs:
                            cpu_0_data_master_granted_row_s1,
                            cpu_0_data_master_qualified_request_row_s1,
                            cpu_0_data_master_read_data_valid_row_s1,
                            cpu_0_data_master_requests_row_s1,
                            d1_row_s1_end_xfer,
                            row_s1_address,
                            row_s1_chipselect,
                            row_s1_readdata_from_sa,
                            row_s1_reset_n,
                            row_s1_write_n,
                            row_s1_writedata
                         )
;

  output           cpu_0_data_master_granted_row_s1;
  output           cpu_0_data_master_qualified_request_row_s1;
  output           cpu_0_data_master_read_data_valid_row_s1;
  output           cpu_0_data_master_requests_row_s1;
  output           d1_row_s1_end_xfer;
  output  [  1: 0] row_s1_address;
  output           row_s1_chipselect;
  output  [ 15: 0] row_s1_readdata_from_sa;
  output           row_s1_reset_n;
  output           row_s1_write_n;
  output  [ 15: 0] row_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input            reset_n;
  input   [ 15: 0] row_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_row_s1;
  wire             cpu_0_data_master_qualified_request_row_s1;
  wire             cpu_0_data_master_read_data_valid_row_s1;
  wire             cpu_0_data_master_requests_row_s1;
  wire             cpu_0_data_master_saved_grant_row_s1;
  reg              d1_reasons_to_wait;
  reg              d1_row_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_row_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  wire    [  1: 0] row_s1_address;
  wire             row_s1_allgrants;
  wire             row_s1_allow_new_arb_cycle;
  wire             row_s1_any_bursting_master_saved_grant;
  wire             row_s1_any_continuerequest;
  wire             row_s1_arb_counter_enable;
  reg     [  1: 0] row_s1_arb_share_counter;
  wire    [  1: 0] row_s1_arb_share_counter_next_value;
  wire    [  1: 0] row_s1_arb_share_set_values;
  wire             row_s1_beginbursttransfer_internal;
  wire             row_s1_begins_xfer;
  wire             row_s1_chipselect;
  wire             row_s1_end_xfer;
  wire             row_s1_firsttransfer;
  wire             row_s1_grant_vector;
  wire             row_s1_in_a_read_cycle;
  wire             row_s1_in_a_write_cycle;
  wire             row_s1_master_qreq_vector;
  wire             row_s1_non_bursting_master_requests;
  wire    [ 15: 0] row_s1_readdata_from_sa;
  reg              row_s1_reg_firsttransfer;
  wire             row_s1_reset_n;
  reg              row_s1_slavearbiterlockenable;
  wire             row_s1_slavearbiterlockenable2;
  wire             row_s1_unreg_firsttransfer;
  wire             row_s1_waits_for_read;
  wire             row_s1_waits_for_write;
  wire             row_s1_write_n;
  wire    [ 15: 0] row_s1_writedata;
  wire    [ 24: 0] shifted_address_to_row_s1_from_cpu_0_data_master;
  wire             wait_for_row_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~row_s1_end_xfer;
    end


  assign row_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_row_s1));
  //assign row_s1_readdata_from_sa = row_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign row_s1_readdata_from_sa = row_s1_readdata;

  assign cpu_0_data_master_requests_row_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010d0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //row_s1_arb_share_counter set values, which is an e_mux
  assign row_s1_arb_share_set_values = 1;

  //row_s1_non_bursting_master_requests mux, which is an e_mux
  assign row_s1_non_bursting_master_requests = cpu_0_data_master_requests_row_s1;

  //row_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign row_s1_any_bursting_master_saved_grant = 0;

  //row_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign row_s1_arb_share_counter_next_value = row_s1_firsttransfer ? (row_s1_arb_share_set_values - 1) : |row_s1_arb_share_counter ? (row_s1_arb_share_counter - 1) : 0;

  //row_s1_allgrants all slave grants, which is an e_mux
  assign row_s1_allgrants = |row_s1_grant_vector;

  //row_s1_end_xfer assignment, which is an e_assign
  assign row_s1_end_xfer = ~(row_s1_waits_for_read | row_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_row_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_row_s1 = row_s1_end_xfer & (~row_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //row_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign row_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_row_s1 & row_s1_allgrants) | (end_xfer_arb_share_counter_term_row_s1 & ~row_s1_non_bursting_master_requests);

  //row_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          row_s1_arb_share_counter <= 0;
      else if (row_s1_arb_counter_enable)
          row_s1_arb_share_counter <= row_s1_arb_share_counter_next_value;
    end


  //row_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          row_s1_slavearbiterlockenable <= 0;
      else if ((|row_s1_master_qreq_vector & end_xfer_arb_share_counter_term_row_s1) | (end_xfer_arb_share_counter_term_row_s1 & ~row_s1_non_bursting_master_requests))
          row_s1_slavearbiterlockenable <= |row_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master row/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = row_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //row_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign row_s1_slavearbiterlockenable2 = |row_s1_arb_share_counter_next_value;

  //cpu_0/data_master row/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = row_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //row_s1_any_continuerequest at least one master continues requesting, which is an e_assign
  assign row_s1_any_continuerequest = 1;

  //cpu_0_data_master_continuerequest continued request, which is an e_assign
  assign cpu_0_data_master_continuerequest = 1;

  assign cpu_0_data_master_qualified_request_row_s1 = cpu_0_data_master_requests_row_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))));
  //local readdatavalid cpu_0_data_master_read_data_valid_row_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_row_s1 = cpu_0_data_master_granted_row_s1 & cpu_0_data_master_read & ~row_s1_waits_for_read;

  //row_s1_writedata mux, which is an e_mux
  assign row_s1_writedata = cpu_0_data_master_writedata;

  //master is always granted when requested
  assign cpu_0_data_master_granted_row_s1 = cpu_0_data_master_qualified_request_row_s1;

  //cpu_0/data_master saved-grant row/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_row_s1 = cpu_0_data_master_requests_row_s1;

  //allow new arb cycle for row/s1, which is an e_assign
  assign row_s1_allow_new_arb_cycle = 1;

  //placeholder chosen master
  assign row_s1_grant_vector = 1;

  //placeholder vector of master qualified-requests
  assign row_s1_master_qreq_vector = 1;

  //row_s1_reset_n assignment, which is an e_assign
  assign row_s1_reset_n = reset_n;

  assign row_s1_chipselect = cpu_0_data_master_granted_row_s1;
  //row_s1_firsttransfer first transaction, which is an e_assign
  assign row_s1_firsttransfer = row_s1_begins_xfer ? row_s1_unreg_firsttransfer : row_s1_reg_firsttransfer;

  //row_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign row_s1_unreg_firsttransfer = ~(row_s1_slavearbiterlockenable & row_s1_any_continuerequest);

  //row_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          row_s1_reg_firsttransfer <= 1'b1;
      else if (row_s1_begins_xfer)
          row_s1_reg_firsttransfer <= row_s1_unreg_firsttransfer;
    end


  //row_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign row_s1_beginbursttransfer_internal = row_s1_begins_xfer;

  //~row_s1_write_n assignment, which is an e_mux
  assign row_s1_write_n = ~(cpu_0_data_master_granted_row_s1 & cpu_0_data_master_write);

  assign shifted_address_to_row_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //row_s1_address mux, which is an e_mux
  assign row_s1_address = shifted_address_to_row_s1_from_cpu_0_data_master >> 2;

  //d1_row_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_row_s1_end_xfer <= 1;
      else 
        d1_row_s1_end_xfer <= row_s1_end_xfer;
    end


  //row_s1_waits_for_read in a cycle, which is an e_mux
  assign row_s1_waits_for_read = row_s1_in_a_read_cycle & row_s1_begins_xfer;

  //row_s1_in_a_read_cycle assignment, which is an e_assign
  assign row_s1_in_a_read_cycle = cpu_0_data_master_granted_row_s1 & cpu_0_data_master_read;

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = row_s1_in_a_read_cycle;

  //row_s1_waits_for_write in a cycle, which is an e_mux
  assign row_s1_waits_for_write = row_s1_in_a_write_cycle & 0;

  //row_s1_in_a_write_cycle assignment, which is an e_assign
  assign row_s1_in_a_write_cycle = cpu_0_data_master_granted_row_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = row_s1_in_a_write_cycle;

  assign wait_for_row_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //row/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_0_data_master_to_sdram_0_s1_module (
                                                             // inputs:
                                                              clear_fifo,
                                                              clk,
                                                              data_in,
                                                              read,
                                                              reset_n,
                                                              sync_reset,
                                                              write,

                                                             // outputs:
                                                              data_out,
                                                              empty,
                                                              fifo_contains_ones_n,
                                                              full
                                                           )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module rdv_fifo_for_cpu_0_instruction_master_to_sdram_0_s1_module (
                                                                    // inputs:
                                                                     clear_fifo,
                                                                     clk,
                                                                     data_in,
                                                                     read,
                                                                     reset_n,
                                                                     sync_reset,
                                                                     write,

                                                                    // outputs:
                                                                     data_out,
                                                                     empty,
                                                                     fifo_contains_ones_n,
                                                                     full
                                                                  )
;

  output           data_out;
  output           empty;
  output           fifo_contains_ones_n;
  output           full;
  input            clear_fifo;
  input            clk;
  input            data_in;
  input            read;
  input            reset_n;
  input            sync_reset;
  input            write;

  wire             data_out;
  wire             empty;
  reg              fifo_contains_ones_n;
  wire             full;
  reg              full_0;
  reg              full_1;
  reg              full_2;
  reg              full_3;
  reg              full_4;
  reg              full_5;
  reg              full_6;
  wire             full_7;
  reg     [  3: 0] how_many_ones;
  wire    [  3: 0] one_count_minus_one;
  wire    [  3: 0] one_count_plus_one;
  wire             p0_full_0;
  wire             p0_stage_0;
  wire             p1_full_1;
  wire             p1_stage_1;
  wire             p2_full_2;
  wire             p2_stage_2;
  wire             p3_full_3;
  wire             p3_stage_3;
  wire             p4_full_4;
  wire             p4_stage_4;
  wire             p5_full_5;
  wire             p5_stage_5;
  wire             p6_full_6;
  wire             p6_stage_6;
  reg              stage_0;
  reg              stage_1;
  reg              stage_2;
  reg              stage_3;
  reg              stage_4;
  reg              stage_5;
  reg              stage_6;
  wire    [  3: 0] updated_one_count;
  assign data_out = stage_0;
  assign full = full_6;
  assign empty = !full_0;
  assign full_7 = 0;
  //data_6, which is an e_mux
  assign p6_stage_6 = ((full_7 & ~clear_fifo) == 0)? data_in :
    data_in;

  //data_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_6 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_6))
          if (sync_reset & full_6 & !((full_7 == 0) & read & write))
              stage_6 <= 0;
          else 
            stage_6 <= p6_stage_6;
    end


  //control_6, which is an e_mux
  assign p6_full_6 = ((read & !write) == 0)? full_5 :
    0;

  //control_reg_6, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_6 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_6 <= 0;
          else 
            full_6 <= p6_full_6;
    end


  //data_5, which is an e_mux
  assign p5_stage_5 = ((full_6 & ~clear_fifo) == 0)? data_in :
    stage_6;

  //data_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_5 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_5))
          if (sync_reset & full_5 & !((full_6 == 0) & read & write))
              stage_5 <= 0;
          else 
            stage_5 <= p5_stage_5;
    end


  //control_5, which is an e_mux
  assign p5_full_5 = ((read & !write) == 0)? full_4 :
    full_6;

  //control_reg_5, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_5 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_5 <= 0;
          else 
            full_5 <= p5_full_5;
    end


  //data_4, which is an e_mux
  assign p4_stage_4 = ((full_5 & ~clear_fifo) == 0)? data_in :
    stage_5;

  //data_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_4 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_4))
          if (sync_reset & full_4 & !((full_5 == 0) & read & write))
              stage_4 <= 0;
          else 
            stage_4 <= p4_stage_4;
    end


  //control_4, which is an e_mux
  assign p4_full_4 = ((read & !write) == 0)? full_3 :
    full_5;

  //control_reg_4, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_4 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_4 <= 0;
          else 
            full_4 <= p4_full_4;
    end


  //data_3, which is an e_mux
  assign p3_stage_3 = ((full_4 & ~clear_fifo) == 0)? data_in :
    stage_4;

  //data_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_3 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_3))
          if (sync_reset & full_3 & !((full_4 == 0) & read & write))
              stage_3 <= 0;
          else 
            stage_3 <= p3_stage_3;
    end


  //control_3, which is an e_mux
  assign p3_full_3 = ((read & !write) == 0)? full_2 :
    full_4;

  //control_reg_3, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_3 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_3 <= 0;
          else 
            full_3 <= p3_full_3;
    end


  //data_2, which is an e_mux
  assign p2_stage_2 = ((full_3 & ~clear_fifo) == 0)? data_in :
    stage_3;

  //data_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_2 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_2))
          if (sync_reset & full_2 & !((full_3 == 0) & read & write))
              stage_2 <= 0;
          else 
            stage_2 <= p2_stage_2;
    end


  //control_2, which is an e_mux
  assign p2_full_2 = ((read & !write) == 0)? full_1 :
    full_3;

  //control_reg_2, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_2 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_2 <= 0;
          else 
            full_2 <= p2_full_2;
    end


  //data_1, which is an e_mux
  assign p1_stage_1 = ((full_2 & ~clear_fifo) == 0)? data_in :
    stage_2;

  //data_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_1 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_1))
          if (sync_reset & full_1 & !((full_2 == 0) & read & write))
              stage_1 <= 0;
          else 
            stage_1 <= p1_stage_1;
    end


  //control_1, which is an e_mux
  assign p1_full_1 = ((read & !write) == 0)? full_0 :
    full_2;

  //control_reg_1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_1 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo)
              full_1 <= 0;
          else 
            full_1 <= p1_full_1;
    end


  //data_0, which is an e_mux
  assign p0_stage_0 = ((full_1 & ~clear_fifo) == 0)? data_in :
    stage_1;

  //data_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          stage_0 <= 0;
      else if (clear_fifo | sync_reset | read | (write & !full_0))
          if (sync_reset & full_0 & !((full_1 == 0) & read & write))
              stage_0 <= 0;
          else 
            stage_0 <= p0_stage_0;
    end


  //control_0, which is an e_mux
  assign p0_full_0 = ((read & !write) == 0)? 1 :
    full_1;

  //control_reg_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          full_0 <= 0;
      else if (clear_fifo | (read ^ write) | (write & !full_0))
          if (clear_fifo & ~write)
              full_0 <= 0;
          else 
            full_0 <= p0_full_0;
    end


  assign one_count_plus_one = how_many_ones + 1;
  assign one_count_minus_one = how_many_ones - 1;
  //updated_one_count, which is an e_mux
  assign updated_one_count = ((((clear_fifo | sync_reset) & !write)))? 0 :
    ((((clear_fifo | sync_reset) & write)))? |data_in :
    ((read & (|data_in) & write & (|stage_0)))? how_many_ones :
    ((write & (|data_in)))? one_count_plus_one :
    ((read & (|stage_0)))? one_count_minus_one :
    how_many_ones;

  //counts how many ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          how_many_ones <= 0;
      else if (clear_fifo | sync_reset | read | write)
          how_many_ones <= updated_one_count;
    end


  //this fifo contains ones in the data pipeline, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          fifo_contains_ones_n <= 1;
      else if (clear_fifo | sync_reset | read | write)
          fifo_contains_ones_n <= ~(|updated_one_count);
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module sdram_0_s1_arbitrator (
                               // inputs:
                                clk,
                                cpu_0_data_master_address_to_slave,
                                cpu_0_data_master_byteenable,
                                cpu_0_data_master_dbs_address,
                                cpu_0_data_master_dbs_write_16,
                                cpu_0_data_master_latency_counter,
                                cpu_0_data_master_read,
                                cpu_0_data_master_write,
                                cpu_0_instruction_master_address_to_slave,
                                cpu_0_instruction_master_dbs_address,
                                cpu_0_instruction_master_latency_counter,
                                cpu_0_instruction_master_read,
                                reset_n,
                                sdram_0_s1_readdata,
                                sdram_0_s1_readdatavalid,
                                sdram_0_s1_waitrequest,

                               // outputs:
                                cpu_0_data_master_byteenable_sdram_0_s1,
                                cpu_0_data_master_granted_sdram_0_s1,
                                cpu_0_data_master_qualified_request_sdram_0_s1,
                                cpu_0_data_master_read_data_valid_sdram_0_s1,
                                cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                cpu_0_data_master_requests_sdram_0_s1,
                                cpu_0_instruction_master_granted_sdram_0_s1,
                                cpu_0_instruction_master_qualified_request_sdram_0_s1,
                                cpu_0_instruction_master_read_data_valid_sdram_0_s1,
                                cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                cpu_0_instruction_master_requests_sdram_0_s1,
                                d1_sdram_0_s1_end_xfer,
                                sdram_0_s1_address,
                                sdram_0_s1_byteenable_n,
                                sdram_0_s1_chipselect,
                                sdram_0_s1_read_n,
                                sdram_0_s1_readdata_from_sa,
                                sdram_0_s1_reset_n,
                                sdram_0_s1_waitrequest_from_sa,
                                sdram_0_s1_write_n,
                                sdram_0_s1_writedata
                             )
;

  output  [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1;
  output           cpu_0_data_master_granted_sdram_0_s1;
  output           cpu_0_data_master_qualified_request_sdram_0_s1;
  output           cpu_0_data_master_read_data_valid_sdram_0_s1;
  output           cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  output           cpu_0_data_master_requests_sdram_0_s1;
  output           cpu_0_instruction_master_granted_sdram_0_s1;
  output           cpu_0_instruction_master_qualified_request_sdram_0_s1;
  output           cpu_0_instruction_master_read_data_valid_sdram_0_s1;
  output           cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  output           cpu_0_instruction_master_requests_sdram_0_s1;
  output           d1_sdram_0_s1_end_xfer;
  output  [ 21: 0] sdram_0_s1_address;
  output  [  1: 0] sdram_0_s1_byteenable_n;
  output           sdram_0_s1_chipselect;
  output           sdram_0_s1_read_n;
  output  [ 15: 0] sdram_0_s1_readdata_from_sa;
  output           sdram_0_s1_reset_n;
  output           sdram_0_s1_waitrequest_from_sa;
  output           sdram_0_s1_write_n;
  output  [ 15: 0] sdram_0_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_dbs_address;
  input   [ 15: 0] cpu_0_data_master_dbs_write_16;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_write;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_dbs_address;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            reset_n;
  input   [ 15: 0] sdram_0_s1_readdata;
  input            sdram_0_s1_readdatavalid;
  input            sdram_0_s1_waitrequest;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire    [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1;
  wire    [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1_segment_0;
  wire    [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1_segment_1;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_sdram_0_s1;
  wire             cpu_0_data_master_qualified_request_sdram_0_s1;
  wire             cpu_0_data_master_rdv_fifo_empty_sdram_0_s1;
  wire             cpu_0_data_master_rdv_fifo_output_from_sdram_0_s1;
  wire             cpu_0_data_master_read_data_valid_sdram_0_s1;
  wire             cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  wire             cpu_0_data_master_requests_sdram_0_s1;
  wire             cpu_0_data_master_saved_grant_sdram_0_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_sdram_0_s1;
  wire             cpu_0_instruction_master_qualified_request_sdram_0_s1;
  wire             cpu_0_instruction_master_rdv_fifo_empty_sdram_0_s1;
  wire             cpu_0_instruction_master_rdv_fifo_output_from_sdram_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_sdram_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  wire             cpu_0_instruction_master_requests_sdram_0_s1;
  wire             cpu_0_instruction_master_saved_grant_sdram_0_s1;
  reg              d1_reasons_to_wait;
  reg              d1_sdram_0_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_sdram_0_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_sdram_0_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_sdram_0_s1;
  wire    [ 21: 0] sdram_0_s1_address;
  wire             sdram_0_s1_allgrants;
  wire             sdram_0_s1_allow_new_arb_cycle;
  wire             sdram_0_s1_any_bursting_master_saved_grant;
  wire             sdram_0_s1_any_continuerequest;
  reg     [  1: 0] sdram_0_s1_arb_addend;
  wire             sdram_0_s1_arb_counter_enable;
  reg     [  1: 0] sdram_0_s1_arb_share_counter;
  wire    [  1: 0] sdram_0_s1_arb_share_counter_next_value;
  wire    [  1: 0] sdram_0_s1_arb_share_set_values;
  wire    [  1: 0] sdram_0_s1_arb_winner;
  wire             sdram_0_s1_arbitration_holdoff_internal;
  wire             sdram_0_s1_beginbursttransfer_internal;
  wire             sdram_0_s1_begins_xfer;
  wire    [  1: 0] sdram_0_s1_byteenable_n;
  wire             sdram_0_s1_chipselect;
  wire    [  3: 0] sdram_0_s1_chosen_master_double_vector;
  wire    [  1: 0] sdram_0_s1_chosen_master_rot_left;
  wire             sdram_0_s1_end_xfer;
  wire             sdram_0_s1_firsttransfer;
  wire    [  1: 0] sdram_0_s1_grant_vector;
  wire             sdram_0_s1_in_a_read_cycle;
  wire             sdram_0_s1_in_a_write_cycle;
  wire    [  1: 0] sdram_0_s1_master_qreq_vector;
  wire             sdram_0_s1_move_on_to_next_transaction;
  wire             sdram_0_s1_non_bursting_master_requests;
  wire             sdram_0_s1_read_n;
  wire    [ 15: 0] sdram_0_s1_readdata_from_sa;
  wire             sdram_0_s1_readdatavalid_from_sa;
  reg              sdram_0_s1_reg_firsttransfer;
  wire             sdram_0_s1_reset_n;
  reg     [  1: 0] sdram_0_s1_saved_chosen_master_vector;
  reg              sdram_0_s1_slavearbiterlockenable;
  wire             sdram_0_s1_slavearbiterlockenable2;
  wire             sdram_0_s1_unreg_firsttransfer;
  wire             sdram_0_s1_waitrequest_from_sa;
  wire             sdram_0_s1_waits_for_read;
  wire             sdram_0_s1_waits_for_write;
  wire             sdram_0_s1_write_n;
  wire    [ 15: 0] sdram_0_s1_writedata;
  wire    [ 24: 0] shifted_address_to_sdram_0_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_sdram_0_s1_from_cpu_0_instruction_master;
  wire             wait_for_sdram_0_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~sdram_0_s1_end_xfer;
    end


  assign sdram_0_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_sdram_0_s1 | cpu_0_instruction_master_qualified_request_sdram_0_s1));
  //assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_readdatavalid_from_sa = sdram_0_s1_readdatavalid;

  //assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_readdata_from_sa = sdram_0_s1_readdata;

  assign cpu_0_data_master_requests_sdram_0_s1 = ({cpu_0_data_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign sdram_0_s1_waitrequest_from_sa = sdram_0_s1_waitrequest;

  //sdram_0_s1_arb_share_counter set values, which is an e_mux
  assign sdram_0_s1_arb_share_set_values = (cpu_0_data_master_granted_sdram_0_s1)? 2 :
    (cpu_0_instruction_master_granted_sdram_0_s1)? 2 :
    (cpu_0_data_master_granted_sdram_0_s1)? 2 :
    (cpu_0_instruction_master_granted_sdram_0_s1)? 2 :
    1;

  //sdram_0_s1_non_bursting_master_requests mux, which is an e_mux
  assign sdram_0_s1_non_bursting_master_requests = cpu_0_data_master_requests_sdram_0_s1 |
    cpu_0_instruction_master_requests_sdram_0_s1 |
    cpu_0_data_master_requests_sdram_0_s1 |
    cpu_0_instruction_master_requests_sdram_0_s1;

  //sdram_0_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign sdram_0_s1_any_bursting_master_saved_grant = 0;

  //sdram_0_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign sdram_0_s1_arb_share_counter_next_value = sdram_0_s1_firsttransfer ? (sdram_0_s1_arb_share_set_values - 1) : |sdram_0_s1_arb_share_counter ? (sdram_0_s1_arb_share_counter - 1) : 0;

  //sdram_0_s1_allgrants all slave grants, which is an e_mux
  assign sdram_0_s1_allgrants = (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector) |
    (|sdram_0_s1_grant_vector);

  //sdram_0_s1_end_xfer assignment, which is an e_assign
  assign sdram_0_s1_end_xfer = ~(sdram_0_s1_waits_for_read | sdram_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_sdram_0_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_sdram_0_s1 = sdram_0_s1_end_xfer & (~sdram_0_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //sdram_0_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign sdram_0_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_sdram_0_s1 & sdram_0_s1_allgrants) | (end_xfer_arb_share_counter_term_sdram_0_s1 & ~sdram_0_s1_non_bursting_master_requests);

  //sdram_0_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_arb_share_counter <= 0;
      else if (sdram_0_s1_arb_counter_enable)
          sdram_0_s1_arb_share_counter <= sdram_0_s1_arb_share_counter_next_value;
    end


  //sdram_0_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_slavearbiterlockenable <= 0;
      else if ((|sdram_0_s1_master_qreq_vector & end_xfer_arb_share_counter_term_sdram_0_s1) | (end_xfer_arb_share_counter_term_sdram_0_s1 & ~sdram_0_s1_non_bursting_master_requests))
          sdram_0_s1_slavearbiterlockenable <= |sdram_0_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master sdram_0/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = sdram_0_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //sdram_0_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign sdram_0_s1_slavearbiterlockenable2 = |sdram_0_s1_arb_share_counter_next_value;

  //cpu_0/data_master sdram_0/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master sdram_0/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = sdram_0_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master sdram_0/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = sdram_0_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_sdram_0_s1 <= cpu_0_instruction_master_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_sdram_0_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_sdram_0_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_sdram_0_s1 & cpu_0_instruction_master_requests_sdram_0_s1;

  //sdram_0_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign sdram_0_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_sdram_0_s1 = cpu_0_data_master_requests_sdram_0_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (1 < cpu_0_data_master_latency_counter))) | ((!cpu_0_data_master_byteenable_sdram_0_s1) & cpu_0_data_master_write) | cpu_0_instruction_master_arbiterlock);
  //unique name for sdram_0_s1_move_on_to_next_transaction, which is an e_assign
  assign sdram_0_s1_move_on_to_next_transaction = sdram_0_s1_readdatavalid_from_sa;

  //rdv_fifo_for_cpu_0_data_master_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_data_master_to_sdram_0_s1_module rdv_fifo_for_cpu_0_data_master_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_0_data_master_granted_sdram_0_s1),
      .data_out             (cpu_0_data_master_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_0_data_master_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register = ~cpu_0_data_master_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid cpu_0_data_master_read_data_valid_sdram_0_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & cpu_0_data_master_rdv_fifo_output_from_sdram_0_s1) & ~ cpu_0_data_master_rdv_fifo_empty_sdram_0_s1;

  //sdram_0_s1_writedata mux, which is an e_mux
  assign sdram_0_s1_writedata = cpu_0_data_master_dbs_write_16;

  assign cpu_0_instruction_master_requests_sdram_0_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 23] , 23'b0} == 25'h800000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted sdram_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_sdram_0_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_sdram_0_s1 <= cpu_0_data_master_saved_grant_sdram_0_s1 ? 1 : (sdram_0_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_sdram_0_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_sdram_0_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_sdram_0_s1 & cpu_0_data_master_requests_sdram_0_s1;

  assign cpu_0_instruction_master_qualified_request_sdram_0_s1 = cpu_0_instruction_master_requests_sdram_0_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (1 < cpu_0_instruction_master_latency_counter))) | cpu_0_data_master_arbiterlock);
  //rdv_fifo_for_cpu_0_instruction_master_to_sdram_0_s1, which is an e_fifo_with_registered_outputs
  rdv_fifo_for_cpu_0_instruction_master_to_sdram_0_s1_module rdv_fifo_for_cpu_0_instruction_master_to_sdram_0_s1
    (
      .clear_fifo           (1'b0),
      .clk                  (clk),
      .data_in              (cpu_0_instruction_master_granted_sdram_0_s1),
      .data_out             (cpu_0_instruction_master_rdv_fifo_output_from_sdram_0_s1),
      .empty                (),
      .fifo_contains_ones_n (cpu_0_instruction_master_rdv_fifo_empty_sdram_0_s1),
      .full                 (),
      .read                 (sdram_0_s1_move_on_to_next_transaction),
      .reset_n              (reset_n),
      .sync_reset           (1'b0),
      .write                (in_a_read_cycle & ~sdram_0_s1_waits_for_read)
    );

  assign cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register = ~cpu_0_instruction_master_rdv_fifo_empty_sdram_0_s1;
  //local readdatavalid cpu_0_instruction_master_read_data_valid_sdram_0_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_sdram_0_s1 = (sdram_0_s1_readdatavalid_from_sa & cpu_0_instruction_master_rdv_fifo_output_from_sdram_0_s1) & ~ cpu_0_instruction_master_rdv_fifo_empty_sdram_0_s1;

  //allow new arb cycle for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_sdram_0_s1;

  //cpu_0/instruction_master grant sdram_0/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_sdram_0_s1 = sdram_0_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant sdram_0/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[0] && cpu_0_instruction_master_requests_sdram_0_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for sdram_0/s1, which is an e_assign
  assign sdram_0_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_sdram_0_s1;

  //cpu_0/data_master grant sdram_0/s1, which is an e_assign
  assign cpu_0_data_master_granted_sdram_0_s1 = sdram_0_s1_grant_vector[1];

  //cpu_0/data_master saved-grant sdram_0/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_sdram_0_s1 = sdram_0_s1_arb_winner[1] && cpu_0_data_master_requests_sdram_0_s1;

  //sdram_0/s1 chosen-master double-vector, which is an e_assign
  assign sdram_0_s1_chosen_master_double_vector = {sdram_0_s1_master_qreq_vector, sdram_0_s1_master_qreq_vector} & ({~sdram_0_s1_master_qreq_vector, ~sdram_0_s1_master_qreq_vector} + sdram_0_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign sdram_0_s1_arb_winner = (sdram_0_s1_allow_new_arb_cycle & | sdram_0_s1_grant_vector) ? sdram_0_s1_grant_vector : sdram_0_s1_saved_chosen_master_vector;

  //saved sdram_0_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_saved_chosen_master_vector <= 0;
      else if (sdram_0_s1_allow_new_arb_cycle)
          sdram_0_s1_saved_chosen_master_vector <= |sdram_0_s1_grant_vector ? sdram_0_s1_grant_vector : sdram_0_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign sdram_0_s1_grant_vector = {(sdram_0_s1_chosen_master_double_vector[1] | sdram_0_s1_chosen_master_double_vector[3]),
    (sdram_0_s1_chosen_master_double_vector[0] | sdram_0_s1_chosen_master_double_vector[2])};

  //sdram_0/s1 chosen master rotated left, which is an e_assign
  assign sdram_0_s1_chosen_master_rot_left = (sdram_0_s1_arb_winner << 1) ? (sdram_0_s1_arb_winner << 1) : 1;

  //sdram_0/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_arb_addend <= 1;
      else if (|sdram_0_s1_grant_vector)
          sdram_0_s1_arb_addend <= sdram_0_s1_end_xfer? sdram_0_s1_chosen_master_rot_left : sdram_0_s1_grant_vector;
    end


  //sdram_0_s1_reset_n assignment, which is an e_assign
  assign sdram_0_s1_reset_n = reset_n;

  assign sdram_0_s1_chipselect = cpu_0_data_master_granted_sdram_0_s1 | cpu_0_instruction_master_granted_sdram_0_s1;
  //sdram_0_s1_firsttransfer first transaction, which is an e_assign
  assign sdram_0_s1_firsttransfer = sdram_0_s1_begins_xfer ? sdram_0_s1_unreg_firsttransfer : sdram_0_s1_reg_firsttransfer;

  //sdram_0_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign sdram_0_s1_unreg_firsttransfer = ~(sdram_0_s1_slavearbiterlockenable & sdram_0_s1_any_continuerequest);

  //sdram_0_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          sdram_0_s1_reg_firsttransfer <= 1'b1;
      else if (sdram_0_s1_begins_xfer)
          sdram_0_s1_reg_firsttransfer <= sdram_0_s1_unreg_firsttransfer;
    end


  //sdram_0_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign sdram_0_s1_beginbursttransfer_internal = sdram_0_s1_begins_xfer;

  //sdram_0_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign sdram_0_s1_arbitration_holdoff_internal = sdram_0_s1_begins_xfer & sdram_0_s1_firsttransfer;

  //~sdram_0_s1_read_n assignment, which is an e_mux
  assign sdram_0_s1_read_n = ~((cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_sdram_0_s1 & cpu_0_instruction_master_read));

  //~sdram_0_s1_write_n assignment, which is an e_mux
  assign sdram_0_s1_write_n = ~(cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_write);

  assign shifted_address_to_sdram_0_s1_from_cpu_0_data_master = {cpu_0_data_master_address_to_slave >> 2,
    cpu_0_data_master_dbs_address[1],
    {1 {1'b0}}};

  //sdram_0_s1_address mux, which is an e_mux
  assign sdram_0_s1_address = (cpu_0_data_master_granted_sdram_0_s1)? (shifted_address_to_sdram_0_s1_from_cpu_0_data_master >> 1) :
    (shifted_address_to_sdram_0_s1_from_cpu_0_instruction_master >> 1);

  assign shifted_address_to_sdram_0_s1_from_cpu_0_instruction_master = {cpu_0_instruction_master_address_to_slave >> 2,
    cpu_0_instruction_master_dbs_address[1],
    {1 {1'b0}}};

  //d1_sdram_0_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_sdram_0_s1_end_xfer <= 1;
      else 
        d1_sdram_0_s1_end_xfer <= sdram_0_s1_end_xfer;
    end


  //sdram_0_s1_waits_for_read in a cycle, which is an e_mux
  assign sdram_0_s1_waits_for_read = sdram_0_s1_in_a_read_cycle & sdram_0_s1_waitrequest_from_sa;

  //sdram_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign sdram_0_s1_in_a_read_cycle = (cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_sdram_0_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = sdram_0_s1_in_a_read_cycle;

  //sdram_0_s1_waits_for_write in a cycle, which is an e_mux
  assign sdram_0_s1_waits_for_write = sdram_0_s1_in_a_write_cycle & sdram_0_s1_waitrequest_from_sa;

  //sdram_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign sdram_0_s1_in_a_write_cycle = cpu_0_data_master_granted_sdram_0_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = sdram_0_s1_in_a_write_cycle;

  assign wait_for_sdram_0_s1_counter = 0;
  //~sdram_0_s1_byteenable_n byte enable port mux, which is an e_mux
  assign sdram_0_s1_byteenable_n = ~((cpu_0_data_master_granted_sdram_0_s1)? cpu_0_data_master_byteenable_sdram_0_s1 :
    -1);

  assign {cpu_0_data_master_byteenable_sdram_0_s1_segment_1,
cpu_0_data_master_byteenable_sdram_0_s1_segment_0} = cpu_0_data_master_byteenable;
  assign cpu_0_data_master_byteenable_sdram_0_s1 = ((cpu_0_data_master_dbs_address[1] == 0))? cpu_0_data_master_byteenable_sdram_0_s1_segment_0 :
    cpu_0_data_master_byteenable_sdram_0_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //sdram_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_sdram_0_s1 + cpu_0_instruction_master_granted_sdram_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_sdram_0_s1 + cpu_0_instruction_master_saved_grant_sdram_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tft_lcd_data_s1_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_0_data_master_address_to_slave,
                                     cpu_0_data_master_byteenable,
                                     cpu_0_data_master_latency_counter,
                                     cpu_0_data_master_read,
                                     cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                     cpu_0_data_master_write,
                                     cpu_0_data_master_writedata,
                                     cpu_0_instruction_master_address_to_slave,
                                     cpu_0_instruction_master_latency_counter,
                                     cpu_0_instruction_master_read,
                                     cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                     reset_n,
                                     tft_lcd_data_s1_readdata,

                                    // outputs:
                                     cpu_0_data_master_granted_tft_lcd_data_s1,
                                     cpu_0_data_master_qualified_request_tft_lcd_data_s1,
                                     cpu_0_data_master_read_data_valid_tft_lcd_data_s1,
                                     cpu_0_data_master_requests_tft_lcd_data_s1,
                                     cpu_0_instruction_master_granted_tft_lcd_data_s1,
                                     cpu_0_instruction_master_qualified_request_tft_lcd_data_s1,
                                     cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1,
                                     cpu_0_instruction_master_requests_tft_lcd_data_s1,
                                     d1_tft_lcd_data_s1_end_xfer,
                                     tft_lcd_data_s1_address,
                                     tft_lcd_data_s1_chipselect,
                                     tft_lcd_data_s1_readdata_from_sa,
                                     tft_lcd_data_s1_reset_n,
                                     tft_lcd_data_s1_write_n,
                                     tft_lcd_data_s1_writedata
                                  )
;

  output           cpu_0_data_master_granted_tft_lcd_data_s1;
  output           cpu_0_data_master_qualified_request_tft_lcd_data_s1;
  output           cpu_0_data_master_read_data_valid_tft_lcd_data_s1;
  output           cpu_0_data_master_requests_tft_lcd_data_s1;
  output           cpu_0_instruction_master_granted_tft_lcd_data_s1;
  output           cpu_0_instruction_master_qualified_request_tft_lcd_data_s1;
  output           cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1;
  output           cpu_0_instruction_master_requests_tft_lcd_data_s1;
  output           d1_tft_lcd_data_s1_end_xfer;
  output  [  1: 0] tft_lcd_data_s1_address;
  output           tft_lcd_data_s1_chipselect;
  output  [  7: 0] tft_lcd_data_s1_readdata_from_sa;
  output           tft_lcd_data_s1_reset_n;
  output           tft_lcd_data_s1_write_n;
  output  [  7: 0] tft_lcd_data_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;
  input   [  7: 0] tft_lcd_data_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_tft_lcd_data_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_data_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_data_s1;
  wire             cpu_0_data_master_requests_tft_lcd_data_s1;
  wire             cpu_0_data_master_saved_grant_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_saved_grant_tft_lcd_data_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tft_lcd_data_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tft_lcd_data_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_tft_lcd_data_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_data_s1;
  wire    [ 24: 0] shifted_address_to_tft_lcd_data_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_tft_lcd_data_s1_from_cpu_0_instruction_master;
  wire    [  1: 0] tft_lcd_data_s1_address;
  wire             tft_lcd_data_s1_allgrants;
  wire             tft_lcd_data_s1_allow_new_arb_cycle;
  wire             tft_lcd_data_s1_any_bursting_master_saved_grant;
  wire             tft_lcd_data_s1_any_continuerequest;
  reg     [  1: 0] tft_lcd_data_s1_arb_addend;
  wire             tft_lcd_data_s1_arb_counter_enable;
  reg     [  1: 0] tft_lcd_data_s1_arb_share_counter;
  wire    [  1: 0] tft_lcd_data_s1_arb_share_counter_next_value;
  wire    [  1: 0] tft_lcd_data_s1_arb_share_set_values;
  wire    [  1: 0] tft_lcd_data_s1_arb_winner;
  wire             tft_lcd_data_s1_arbitration_holdoff_internal;
  wire             tft_lcd_data_s1_beginbursttransfer_internal;
  wire             tft_lcd_data_s1_begins_xfer;
  wire             tft_lcd_data_s1_chipselect;
  wire    [  3: 0] tft_lcd_data_s1_chosen_master_double_vector;
  wire    [  1: 0] tft_lcd_data_s1_chosen_master_rot_left;
  wire             tft_lcd_data_s1_end_xfer;
  wire             tft_lcd_data_s1_firsttransfer;
  wire    [  1: 0] tft_lcd_data_s1_grant_vector;
  wire             tft_lcd_data_s1_in_a_read_cycle;
  wire             tft_lcd_data_s1_in_a_write_cycle;
  wire    [  1: 0] tft_lcd_data_s1_master_qreq_vector;
  wire             tft_lcd_data_s1_non_bursting_master_requests;
  wire             tft_lcd_data_s1_pretend_byte_enable;
  wire    [  7: 0] tft_lcd_data_s1_readdata_from_sa;
  reg              tft_lcd_data_s1_reg_firsttransfer;
  wire             tft_lcd_data_s1_reset_n;
  reg     [  1: 0] tft_lcd_data_s1_saved_chosen_master_vector;
  reg              tft_lcd_data_s1_slavearbiterlockenable;
  wire             tft_lcd_data_s1_slavearbiterlockenable2;
  wire             tft_lcd_data_s1_unreg_firsttransfer;
  wire             tft_lcd_data_s1_waits_for_read;
  wire             tft_lcd_data_s1_waits_for_write;
  wire             tft_lcd_data_s1_write_n;
  wire    [  7: 0] tft_lcd_data_s1_writedata;
  wire             wait_for_tft_lcd_data_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tft_lcd_data_s1_end_xfer;
    end


  assign tft_lcd_data_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_tft_lcd_data_s1 | cpu_0_instruction_master_qualified_request_tft_lcd_data_s1));
  //assign tft_lcd_data_s1_readdata_from_sa = tft_lcd_data_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tft_lcd_data_s1_readdata_from_sa = tft_lcd_data_s1_readdata;

  assign cpu_0_data_master_requests_tft_lcd_data_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801070) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //tft_lcd_data_s1_arb_share_counter set values, which is an e_mux
  assign tft_lcd_data_s1_arb_share_set_values = 1;

  //tft_lcd_data_s1_non_bursting_master_requests mux, which is an e_mux
  assign tft_lcd_data_s1_non_bursting_master_requests = cpu_0_data_master_requests_tft_lcd_data_s1 |
    cpu_0_instruction_master_requests_tft_lcd_data_s1 |
    cpu_0_data_master_requests_tft_lcd_data_s1 |
    cpu_0_instruction_master_requests_tft_lcd_data_s1;

  //tft_lcd_data_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tft_lcd_data_s1_any_bursting_master_saved_grant = 0;

  //tft_lcd_data_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tft_lcd_data_s1_arb_share_counter_next_value = tft_lcd_data_s1_firsttransfer ? (tft_lcd_data_s1_arb_share_set_values - 1) : |tft_lcd_data_s1_arb_share_counter ? (tft_lcd_data_s1_arb_share_counter - 1) : 0;

  //tft_lcd_data_s1_allgrants all slave grants, which is an e_mux
  assign tft_lcd_data_s1_allgrants = (|tft_lcd_data_s1_grant_vector) |
    (|tft_lcd_data_s1_grant_vector) |
    (|tft_lcd_data_s1_grant_vector) |
    (|tft_lcd_data_s1_grant_vector);

  //tft_lcd_data_s1_end_xfer assignment, which is an e_assign
  assign tft_lcd_data_s1_end_xfer = ~(tft_lcd_data_s1_waits_for_read | tft_lcd_data_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tft_lcd_data_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tft_lcd_data_s1 = tft_lcd_data_s1_end_xfer & (~tft_lcd_data_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tft_lcd_data_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tft_lcd_data_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tft_lcd_data_s1 & tft_lcd_data_s1_allgrants) | (end_xfer_arb_share_counter_term_tft_lcd_data_s1 & ~tft_lcd_data_s1_non_bursting_master_requests);

  //tft_lcd_data_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_data_s1_arb_share_counter <= 0;
      else if (tft_lcd_data_s1_arb_counter_enable)
          tft_lcd_data_s1_arb_share_counter <= tft_lcd_data_s1_arb_share_counter_next_value;
    end


  //tft_lcd_data_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_data_s1_slavearbiterlockenable <= 0;
      else if ((|tft_lcd_data_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tft_lcd_data_s1) | (end_xfer_arb_share_counter_term_tft_lcd_data_s1 & ~tft_lcd_data_s1_non_bursting_master_requests))
          tft_lcd_data_s1_slavearbiterlockenable <= |tft_lcd_data_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master tft_lcd_data/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tft_lcd_data_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tft_lcd_data_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tft_lcd_data_s1_slavearbiterlockenable2 = |tft_lcd_data_s1_arb_share_counter_next_value;

  //cpu_0/data_master tft_lcd_data/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tft_lcd_data_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_data/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tft_lcd_data_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_data/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tft_lcd_data_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted tft_lcd_data/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_data_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_data_s1 <= cpu_0_instruction_master_saved_grant_tft_lcd_data_s1 ? 1 : (tft_lcd_data_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_tft_lcd_data_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_data_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_data_s1 & cpu_0_instruction_master_requests_tft_lcd_data_s1;

  //tft_lcd_data_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tft_lcd_data_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_tft_lcd_data_s1 = cpu_0_data_master_requests_tft_lcd_data_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_tft_lcd_data_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_tft_lcd_data_s1 = cpu_0_data_master_granted_tft_lcd_data_s1 & cpu_0_data_master_read & ~tft_lcd_data_s1_waits_for_read;

  //tft_lcd_data_s1_writedata mux, which is an e_mux
  assign tft_lcd_data_s1_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_tft_lcd_data_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801070) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted tft_lcd_data/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_tft_lcd_data_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_tft_lcd_data_s1 <= cpu_0_data_master_saved_grant_tft_lcd_data_s1 ? 1 : (tft_lcd_data_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_tft_lcd_data_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_tft_lcd_data_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_tft_lcd_data_s1 & cpu_0_data_master_requests_tft_lcd_data_s1;

  assign cpu_0_instruction_master_qualified_request_tft_lcd_data_s1 = cpu_0_instruction_master_requests_tft_lcd_data_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1 = cpu_0_instruction_master_granted_tft_lcd_data_s1 & cpu_0_instruction_master_read & ~tft_lcd_data_s1_waits_for_read;

  //allow new arb cycle for tft_lcd_data/s1, which is an e_assign
  assign tft_lcd_data_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for tft_lcd_data/s1, which is an e_assign
  assign tft_lcd_data_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_tft_lcd_data_s1;

  //cpu_0/instruction_master grant tft_lcd_data/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_tft_lcd_data_s1 = tft_lcd_data_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant tft_lcd_data/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_tft_lcd_data_s1 = tft_lcd_data_s1_arb_winner[0] && cpu_0_instruction_master_requests_tft_lcd_data_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for tft_lcd_data/s1, which is an e_assign
  assign tft_lcd_data_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_tft_lcd_data_s1;

  //cpu_0/data_master grant tft_lcd_data/s1, which is an e_assign
  assign cpu_0_data_master_granted_tft_lcd_data_s1 = tft_lcd_data_s1_grant_vector[1];

  //cpu_0/data_master saved-grant tft_lcd_data/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_tft_lcd_data_s1 = tft_lcd_data_s1_arb_winner[1] && cpu_0_data_master_requests_tft_lcd_data_s1;

  //tft_lcd_data/s1 chosen-master double-vector, which is an e_assign
  assign tft_lcd_data_s1_chosen_master_double_vector = {tft_lcd_data_s1_master_qreq_vector, tft_lcd_data_s1_master_qreq_vector} & ({~tft_lcd_data_s1_master_qreq_vector, ~tft_lcd_data_s1_master_qreq_vector} + tft_lcd_data_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign tft_lcd_data_s1_arb_winner = (tft_lcd_data_s1_allow_new_arb_cycle & | tft_lcd_data_s1_grant_vector) ? tft_lcd_data_s1_grant_vector : tft_lcd_data_s1_saved_chosen_master_vector;

  //saved tft_lcd_data_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_data_s1_saved_chosen_master_vector <= 0;
      else if (tft_lcd_data_s1_allow_new_arb_cycle)
          tft_lcd_data_s1_saved_chosen_master_vector <= |tft_lcd_data_s1_grant_vector ? tft_lcd_data_s1_grant_vector : tft_lcd_data_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tft_lcd_data_s1_grant_vector = {(tft_lcd_data_s1_chosen_master_double_vector[1] | tft_lcd_data_s1_chosen_master_double_vector[3]),
    (tft_lcd_data_s1_chosen_master_double_vector[0] | tft_lcd_data_s1_chosen_master_double_vector[2])};

  //tft_lcd_data/s1 chosen master rotated left, which is an e_assign
  assign tft_lcd_data_s1_chosen_master_rot_left = (tft_lcd_data_s1_arb_winner << 1) ? (tft_lcd_data_s1_arb_winner << 1) : 1;

  //tft_lcd_data/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_data_s1_arb_addend <= 1;
      else if (|tft_lcd_data_s1_grant_vector)
          tft_lcd_data_s1_arb_addend <= tft_lcd_data_s1_end_xfer? tft_lcd_data_s1_chosen_master_rot_left : tft_lcd_data_s1_grant_vector;
    end


  //tft_lcd_data_s1_reset_n assignment, which is an e_assign
  assign tft_lcd_data_s1_reset_n = reset_n;

  assign tft_lcd_data_s1_chipselect = cpu_0_data_master_granted_tft_lcd_data_s1 | cpu_0_instruction_master_granted_tft_lcd_data_s1;
  //tft_lcd_data_s1_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_data_s1_firsttransfer = tft_lcd_data_s1_begins_xfer ? tft_lcd_data_s1_unreg_firsttransfer : tft_lcd_data_s1_reg_firsttransfer;

  //tft_lcd_data_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_data_s1_unreg_firsttransfer = ~(tft_lcd_data_s1_slavearbiterlockenable & tft_lcd_data_s1_any_continuerequest);

  //tft_lcd_data_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_data_s1_reg_firsttransfer <= 1'b1;
      else if (tft_lcd_data_s1_begins_xfer)
          tft_lcd_data_s1_reg_firsttransfer <= tft_lcd_data_s1_unreg_firsttransfer;
    end


  //tft_lcd_data_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tft_lcd_data_s1_beginbursttransfer_internal = tft_lcd_data_s1_begins_xfer;

  //tft_lcd_data_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tft_lcd_data_s1_arbitration_holdoff_internal = tft_lcd_data_s1_begins_xfer & tft_lcd_data_s1_firsttransfer;

  //~tft_lcd_data_s1_write_n assignment, which is an e_mux
  assign tft_lcd_data_s1_write_n = ~(((cpu_0_data_master_granted_tft_lcd_data_s1 & cpu_0_data_master_write)) & tft_lcd_data_s1_pretend_byte_enable);

  assign shifted_address_to_tft_lcd_data_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //tft_lcd_data_s1_address mux, which is an e_mux
  assign tft_lcd_data_s1_address = (cpu_0_data_master_granted_tft_lcd_data_s1)? (shifted_address_to_tft_lcd_data_s1_from_cpu_0_data_master >> 2) :
    (shifted_address_to_tft_lcd_data_s1_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_tft_lcd_data_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_tft_lcd_data_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tft_lcd_data_s1_end_xfer <= 1;
      else 
        d1_tft_lcd_data_s1_end_xfer <= tft_lcd_data_s1_end_xfer;
    end


  //tft_lcd_data_s1_waits_for_read in a cycle, which is an e_mux
  assign tft_lcd_data_s1_waits_for_read = tft_lcd_data_s1_in_a_read_cycle & tft_lcd_data_s1_begins_xfer;

  //tft_lcd_data_s1_in_a_read_cycle assignment, which is an e_assign
  assign tft_lcd_data_s1_in_a_read_cycle = (cpu_0_data_master_granted_tft_lcd_data_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_tft_lcd_data_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tft_lcd_data_s1_in_a_read_cycle;

  //tft_lcd_data_s1_waits_for_write in a cycle, which is an e_mux
  assign tft_lcd_data_s1_waits_for_write = tft_lcd_data_s1_in_a_write_cycle & 0;

  //tft_lcd_data_s1_in_a_write_cycle assignment, which is an e_assign
  assign tft_lcd_data_s1_in_a_write_cycle = cpu_0_data_master_granted_tft_lcd_data_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tft_lcd_data_s1_in_a_write_cycle;

  assign wait_for_tft_lcd_data_s1_counter = 0;
  //tft_lcd_data_s1_pretend_byte_enable byte enable port mux, which is an e_mux
  assign tft_lcd_data_s1_pretend_byte_enable = (cpu_0_data_master_granted_tft_lcd_data_s1)? cpu_0_data_master_byteenable :
    -1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tft_lcd_data/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_tft_lcd_data_s1 + cpu_0_instruction_master_granted_tft_lcd_data_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_tft_lcd_data_s1 + cpu_0_instruction_master_saved_grant_tft_lcd_data_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tft_lcd_nrd_s1_arbitrator (
                                   // inputs:
                                    clk,
                                    cpu_0_data_master_address_to_slave,
                                    cpu_0_data_master_latency_counter,
                                    cpu_0_data_master_read,
                                    cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                    cpu_0_data_master_write,
                                    cpu_0_data_master_writedata,
                                    cpu_0_instruction_master_address_to_slave,
                                    cpu_0_instruction_master_latency_counter,
                                    cpu_0_instruction_master_read,
                                    cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                    reset_n,
                                    tft_lcd_nrd_s1_readdata,

                                   // outputs:
                                    cpu_0_data_master_granted_tft_lcd_nrd_s1,
                                    cpu_0_data_master_qualified_request_tft_lcd_nrd_s1,
                                    cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1,
                                    cpu_0_data_master_requests_tft_lcd_nrd_s1,
                                    cpu_0_instruction_master_granted_tft_lcd_nrd_s1,
                                    cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1,
                                    cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1,
                                    cpu_0_instruction_master_requests_tft_lcd_nrd_s1,
                                    d1_tft_lcd_nrd_s1_end_xfer,
                                    tft_lcd_nrd_s1_address,
                                    tft_lcd_nrd_s1_chipselect,
                                    tft_lcd_nrd_s1_readdata_from_sa,
                                    tft_lcd_nrd_s1_reset_n,
                                    tft_lcd_nrd_s1_write_n,
                                    tft_lcd_nrd_s1_writedata
                                 )
;

  output           cpu_0_data_master_granted_tft_lcd_nrd_s1;
  output           cpu_0_data_master_qualified_request_tft_lcd_nrd_s1;
  output           cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1;
  output           cpu_0_data_master_requests_tft_lcd_nrd_s1;
  output           cpu_0_instruction_master_granted_tft_lcd_nrd_s1;
  output           cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1;
  output           cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1;
  output           cpu_0_instruction_master_requests_tft_lcd_nrd_s1;
  output           d1_tft_lcd_nrd_s1_end_xfer;
  output  [  1: 0] tft_lcd_nrd_s1_address;
  output           tft_lcd_nrd_s1_chipselect;
  output           tft_lcd_nrd_s1_readdata_from_sa;
  output           tft_lcd_nrd_s1_reset_n;
  output           tft_lcd_nrd_s1_write_n;
  output           tft_lcd_nrd_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;
  input            tft_lcd_nrd_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_saved_grant_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_saved_grant_tft_lcd_nrd_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tft_lcd_nrd_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tft_lcd_nrd_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrd_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrd_s1;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_instruction_master;
  wire    [  1: 0] tft_lcd_nrd_s1_address;
  wire             tft_lcd_nrd_s1_allgrants;
  wire             tft_lcd_nrd_s1_allow_new_arb_cycle;
  wire             tft_lcd_nrd_s1_any_bursting_master_saved_grant;
  wire             tft_lcd_nrd_s1_any_continuerequest;
  reg     [  1: 0] tft_lcd_nrd_s1_arb_addend;
  wire             tft_lcd_nrd_s1_arb_counter_enable;
  reg     [  1: 0] tft_lcd_nrd_s1_arb_share_counter;
  wire    [  1: 0] tft_lcd_nrd_s1_arb_share_counter_next_value;
  wire    [  1: 0] tft_lcd_nrd_s1_arb_share_set_values;
  wire    [  1: 0] tft_lcd_nrd_s1_arb_winner;
  wire             tft_lcd_nrd_s1_arbitration_holdoff_internal;
  wire             tft_lcd_nrd_s1_beginbursttransfer_internal;
  wire             tft_lcd_nrd_s1_begins_xfer;
  wire             tft_lcd_nrd_s1_chipselect;
  wire    [  3: 0] tft_lcd_nrd_s1_chosen_master_double_vector;
  wire    [  1: 0] tft_lcd_nrd_s1_chosen_master_rot_left;
  wire             tft_lcd_nrd_s1_end_xfer;
  wire             tft_lcd_nrd_s1_firsttransfer;
  wire    [  1: 0] tft_lcd_nrd_s1_grant_vector;
  wire             tft_lcd_nrd_s1_in_a_read_cycle;
  wire             tft_lcd_nrd_s1_in_a_write_cycle;
  wire    [  1: 0] tft_lcd_nrd_s1_master_qreq_vector;
  wire             tft_lcd_nrd_s1_non_bursting_master_requests;
  wire             tft_lcd_nrd_s1_readdata_from_sa;
  reg              tft_lcd_nrd_s1_reg_firsttransfer;
  wire             tft_lcd_nrd_s1_reset_n;
  reg     [  1: 0] tft_lcd_nrd_s1_saved_chosen_master_vector;
  reg              tft_lcd_nrd_s1_slavearbiterlockenable;
  wire             tft_lcd_nrd_s1_slavearbiterlockenable2;
  wire             tft_lcd_nrd_s1_unreg_firsttransfer;
  wire             tft_lcd_nrd_s1_waits_for_read;
  wire             tft_lcd_nrd_s1_waits_for_write;
  wire             tft_lcd_nrd_s1_write_n;
  wire             tft_lcd_nrd_s1_writedata;
  wire             wait_for_tft_lcd_nrd_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tft_lcd_nrd_s1_end_xfer;
    end


  assign tft_lcd_nrd_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 | cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1));
  //assign tft_lcd_nrd_s1_readdata_from_sa = tft_lcd_nrd_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tft_lcd_nrd_s1_readdata_from_sa = tft_lcd_nrd_s1_readdata;

  assign cpu_0_data_master_requests_tft_lcd_nrd_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010a0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //tft_lcd_nrd_s1_arb_share_counter set values, which is an e_mux
  assign tft_lcd_nrd_s1_arb_share_set_values = 1;

  //tft_lcd_nrd_s1_non_bursting_master_requests mux, which is an e_mux
  assign tft_lcd_nrd_s1_non_bursting_master_requests = cpu_0_data_master_requests_tft_lcd_nrd_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nrd_s1 |
    cpu_0_data_master_requests_tft_lcd_nrd_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nrd_s1;

  //tft_lcd_nrd_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tft_lcd_nrd_s1_any_bursting_master_saved_grant = 0;

  //tft_lcd_nrd_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tft_lcd_nrd_s1_arb_share_counter_next_value = tft_lcd_nrd_s1_firsttransfer ? (tft_lcd_nrd_s1_arb_share_set_values - 1) : |tft_lcd_nrd_s1_arb_share_counter ? (tft_lcd_nrd_s1_arb_share_counter - 1) : 0;

  //tft_lcd_nrd_s1_allgrants all slave grants, which is an e_mux
  assign tft_lcd_nrd_s1_allgrants = (|tft_lcd_nrd_s1_grant_vector) |
    (|tft_lcd_nrd_s1_grant_vector) |
    (|tft_lcd_nrd_s1_grant_vector) |
    (|tft_lcd_nrd_s1_grant_vector);

  //tft_lcd_nrd_s1_end_xfer assignment, which is an e_assign
  assign tft_lcd_nrd_s1_end_xfer = ~(tft_lcd_nrd_s1_waits_for_read | tft_lcd_nrd_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tft_lcd_nrd_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tft_lcd_nrd_s1 = tft_lcd_nrd_s1_end_xfer & (~tft_lcd_nrd_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tft_lcd_nrd_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tft_lcd_nrd_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tft_lcd_nrd_s1 & tft_lcd_nrd_s1_allgrants) | (end_xfer_arb_share_counter_term_tft_lcd_nrd_s1 & ~tft_lcd_nrd_s1_non_bursting_master_requests);

  //tft_lcd_nrd_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrd_s1_arb_share_counter <= 0;
      else if (tft_lcd_nrd_s1_arb_counter_enable)
          tft_lcd_nrd_s1_arb_share_counter <= tft_lcd_nrd_s1_arb_share_counter_next_value;
    end


  //tft_lcd_nrd_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrd_s1_slavearbiterlockenable <= 0;
      else if ((|tft_lcd_nrd_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tft_lcd_nrd_s1) | (end_xfer_arb_share_counter_term_tft_lcd_nrd_s1 & ~tft_lcd_nrd_s1_non_bursting_master_requests))
          tft_lcd_nrd_s1_slavearbiterlockenable <= |tft_lcd_nrd_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master tft_lcd_nrd/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tft_lcd_nrd_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tft_lcd_nrd_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tft_lcd_nrd_s1_slavearbiterlockenable2 = |tft_lcd_nrd_s1_arb_share_counter_next_value;

  //cpu_0/data_master tft_lcd_nrd/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tft_lcd_nrd_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nrd/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tft_lcd_nrd_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nrd/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tft_lcd_nrd_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted tft_lcd_nrd/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrd_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrd_s1 <= cpu_0_instruction_master_saved_grant_tft_lcd_nrd_s1 ? 1 : (tft_lcd_nrd_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_tft_lcd_nrd_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrd_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrd_s1 & cpu_0_instruction_master_requests_tft_lcd_nrd_s1;

  //tft_lcd_nrd_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tft_lcd_nrd_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_tft_lcd_nrd_s1 = cpu_0_data_master_requests_tft_lcd_nrd_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1 = cpu_0_data_master_granted_tft_lcd_nrd_s1 & cpu_0_data_master_read & ~tft_lcd_nrd_s1_waits_for_read;

  //tft_lcd_nrd_s1_writedata mux, which is an e_mux
  assign tft_lcd_nrd_s1_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_tft_lcd_nrd_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010a0) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted tft_lcd_nrd/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrd_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrd_s1 <= cpu_0_data_master_saved_grant_tft_lcd_nrd_s1 ? 1 : (tft_lcd_nrd_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_tft_lcd_nrd_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrd_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrd_s1 & cpu_0_data_master_requests_tft_lcd_nrd_s1;

  assign cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1 = cpu_0_instruction_master_requests_tft_lcd_nrd_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1 = cpu_0_instruction_master_granted_tft_lcd_nrd_s1 & cpu_0_instruction_master_read & ~tft_lcd_nrd_s1_waits_for_read;

  //allow new arb cycle for tft_lcd_nrd/s1, which is an e_assign
  assign tft_lcd_nrd_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for tft_lcd_nrd/s1, which is an e_assign
  assign tft_lcd_nrd_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1;

  //cpu_0/instruction_master grant tft_lcd_nrd/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_tft_lcd_nrd_s1 = tft_lcd_nrd_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant tft_lcd_nrd/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_tft_lcd_nrd_s1 = tft_lcd_nrd_s1_arb_winner[0] && cpu_0_instruction_master_requests_tft_lcd_nrd_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for tft_lcd_nrd/s1, which is an e_assign
  assign tft_lcd_nrd_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_tft_lcd_nrd_s1;

  //cpu_0/data_master grant tft_lcd_nrd/s1, which is an e_assign
  assign cpu_0_data_master_granted_tft_lcd_nrd_s1 = tft_lcd_nrd_s1_grant_vector[1];

  //cpu_0/data_master saved-grant tft_lcd_nrd/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_tft_lcd_nrd_s1 = tft_lcd_nrd_s1_arb_winner[1] && cpu_0_data_master_requests_tft_lcd_nrd_s1;

  //tft_lcd_nrd/s1 chosen-master double-vector, which is an e_assign
  assign tft_lcd_nrd_s1_chosen_master_double_vector = {tft_lcd_nrd_s1_master_qreq_vector, tft_lcd_nrd_s1_master_qreq_vector} & ({~tft_lcd_nrd_s1_master_qreq_vector, ~tft_lcd_nrd_s1_master_qreq_vector} + tft_lcd_nrd_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign tft_lcd_nrd_s1_arb_winner = (tft_lcd_nrd_s1_allow_new_arb_cycle & | tft_lcd_nrd_s1_grant_vector) ? tft_lcd_nrd_s1_grant_vector : tft_lcd_nrd_s1_saved_chosen_master_vector;

  //saved tft_lcd_nrd_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrd_s1_saved_chosen_master_vector <= 0;
      else if (tft_lcd_nrd_s1_allow_new_arb_cycle)
          tft_lcd_nrd_s1_saved_chosen_master_vector <= |tft_lcd_nrd_s1_grant_vector ? tft_lcd_nrd_s1_grant_vector : tft_lcd_nrd_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tft_lcd_nrd_s1_grant_vector = {(tft_lcd_nrd_s1_chosen_master_double_vector[1] | tft_lcd_nrd_s1_chosen_master_double_vector[3]),
    (tft_lcd_nrd_s1_chosen_master_double_vector[0] | tft_lcd_nrd_s1_chosen_master_double_vector[2])};

  //tft_lcd_nrd/s1 chosen master rotated left, which is an e_assign
  assign tft_lcd_nrd_s1_chosen_master_rot_left = (tft_lcd_nrd_s1_arb_winner << 1) ? (tft_lcd_nrd_s1_arb_winner << 1) : 1;

  //tft_lcd_nrd/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrd_s1_arb_addend <= 1;
      else if (|tft_lcd_nrd_s1_grant_vector)
          tft_lcd_nrd_s1_arb_addend <= tft_lcd_nrd_s1_end_xfer? tft_lcd_nrd_s1_chosen_master_rot_left : tft_lcd_nrd_s1_grant_vector;
    end


  //tft_lcd_nrd_s1_reset_n assignment, which is an e_assign
  assign tft_lcd_nrd_s1_reset_n = reset_n;

  assign tft_lcd_nrd_s1_chipselect = cpu_0_data_master_granted_tft_lcd_nrd_s1 | cpu_0_instruction_master_granted_tft_lcd_nrd_s1;
  //tft_lcd_nrd_s1_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nrd_s1_firsttransfer = tft_lcd_nrd_s1_begins_xfer ? tft_lcd_nrd_s1_unreg_firsttransfer : tft_lcd_nrd_s1_reg_firsttransfer;

  //tft_lcd_nrd_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nrd_s1_unreg_firsttransfer = ~(tft_lcd_nrd_s1_slavearbiterlockenable & tft_lcd_nrd_s1_any_continuerequest);

  //tft_lcd_nrd_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrd_s1_reg_firsttransfer <= 1'b1;
      else if (tft_lcd_nrd_s1_begins_xfer)
          tft_lcd_nrd_s1_reg_firsttransfer <= tft_lcd_nrd_s1_unreg_firsttransfer;
    end


  //tft_lcd_nrd_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tft_lcd_nrd_s1_beginbursttransfer_internal = tft_lcd_nrd_s1_begins_xfer;

  //tft_lcd_nrd_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tft_lcd_nrd_s1_arbitration_holdoff_internal = tft_lcd_nrd_s1_begins_xfer & tft_lcd_nrd_s1_firsttransfer;

  //~tft_lcd_nrd_s1_write_n assignment, which is an e_mux
  assign tft_lcd_nrd_s1_write_n = ~(cpu_0_data_master_granted_tft_lcd_nrd_s1 & cpu_0_data_master_write);

  assign shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //tft_lcd_nrd_s1_address mux, which is an e_mux
  assign tft_lcd_nrd_s1_address = (cpu_0_data_master_granted_tft_lcd_nrd_s1)? (shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_data_master >> 2) :
    (shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_tft_lcd_nrd_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_tft_lcd_nrd_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tft_lcd_nrd_s1_end_xfer <= 1;
      else 
        d1_tft_lcd_nrd_s1_end_xfer <= tft_lcd_nrd_s1_end_xfer;
    end


  //tft_lcd_nrd_s1_waits_for_read in a cycle, which is an e_mux
  assign tft_lcd_nrd_s1_waits_for_read = tft_lcd_nrd_s1_in_a_read_cycle & tft_lcd_nrd_s1_begins_xfer;

  //tft_lcd_nrd_s1_in_a_read_cycle assignment, which is an e_assign
  assign tft_lcd_nrd_s1_in_a_read_cycle = (cpu_0_data_master_granted_tft_lcd_nrd_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_tft_lcd_nrd_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tft_lcd_nrd_s1_in_a_read_cycle;

  //tft_lcd_nrd_s1_waits_for_write in a cycle, which is an e_mux
  assign tft_lcd_nrd_s1_waits_for_write = tft_lcd_nrd_s1_in_a_write_cycle & 0;

  //tft_lcd_nrd_s1_in_a_write_cycle assignment, which is an e_assign
  assign tft_lcd_nrd_s1_in_a_write_cycle = cpu_0_data_master_granted_tft_lcd_nrd_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tft_lcd_nrd_s1_in_a_write_cycle;

  assign wait_for_tft_lcd_nrd_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tft_lcd_nrd/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_tft_lcd_nrd_s1 + cpu_0_instruction_master_granted_tft_lcd_nrd_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_tft_lcd_nrd_s1 + cpu_0_instruction_master_saved_grant_tft_lcd_nrd_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tft_lcd_nrst_s1_arbitrator (
                                    // inputs:
                                     clk,
                                     cpu_0_data_master_address_to_slave,
                                     cpu_0_data_master_latency_counter,
                                     cpu_0_data_master_read,
                                     cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                     cpu_0_data_master_write,
                                     cpu_0_data_master_writedata,
                                     cpu_0_instruction_master_address_to_slave,
                                     cpu_0_instruction_master_latency_counter,
                                     cpu_0_instruction_master_read,
                                     cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                     reset_n,
                                     tft_lcd_nrst_s1_readdata,

                                    // outputs:
                                     cpu_0_data_master_granted_tft_lcd_nrst_s1,
                                     cpu_0_data_master_qualified_request_tft_lcd_nrst_s1,
                                     cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1,
                                     cpu_0_data_master_requests_tft_lcd_nrst_s1,
                                     cpu_0_instruction_master_granted_tft_lcd_nrst_s1,
                                     cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1,
                                     cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1,
                                     cpu_0_instruction_master_requests_tft_lcd_nrst_s1,
                                     d1_tft_lcd_nrst_s1_end_xfer,
                                     tft_lcd_nrst_s1_address,
                                     tft_lcd_nrst_s1_chipselect,
                                     tft_lcd_nrst_s1_readdata_from_sa,
                                     tft_lcd_nrst_s1_reset_n,
                                     tft_lcd_nrst_s1_write_n,
                                     tft_lcd_nrst_s1_writedata
                                  )
;

  output           cpu_0_data_master_granted_tft_lcd_nrst_s1;
  output           cpu_0_data_master_qualified_request_tft_lcd_nrst_s1;
  output           cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1;
  output           cpu_0_data_master_requests_tft_lcd_nrst_s1;
  output           cpu_0_instruction_master_granted_tft_lcd_nrst_s1;
  output           cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1;
  output           cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1;
  output           cpu_0_instruction_master_requests_tft_lcd_nrst_s1;
  output           d1_tft_lcd_nrst_s1_end_xfer;
  output  [  1: 0] tft_lcd_nrst_s1_address;
  output           tft_lcd_nrst_s1_chipselect;
  output           tft_lcd_nrst_s1_readdata_from_sa;
  output           tft_lcd_nrst_s1_reset_n;
  output           tft_lcd_nrst_s1_write_n;
  output           tft_lcd_nrst_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;
  input            tft_lcd_nrst_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_saved_grant_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_saved_grant_tft_lcd_nrst_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tft_lcd_nrst_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tft_lcd_nrst_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrst_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrst_s1;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_instruction_master;
  wire    [  1: 0] tft_lcd_nrst_s1_address;
  wire             tft_lcd_nrst_s1_allgrants;
  wire             tft_lcd_nrst_s1_allow_new_arb_cycle;
  wire             tft_lcd_nrst_s1_any_bursting_master_saved_grant;
  wire             tft_lcd_nrst_s1_any_continuerequest;
  reg     [  1: 0] tft_lcd_nrst_s1_arb_addend;
  wire             tft_lcd_nrst_s1_arb_counter_enable;
  reg     [  1: 0] tft_lcd_nrst_s1_arb_share_counter;
  wire    [  1: 0] tft_lcd_nrst_s1_arb_share_counter_next_value;
  wire    [  1: 0] tft_lcd_nrst_s1_arb_share_set_values;
  wire    [  1: 0] tft_lcd_nrst_s1_arb_winner;
  wire             tft_lcd_nrst_s1_arbitration_holdoff_internal;
  wire             tft_lcd_nrst_s1_beginbursttransfer_internal;
  wire             tft_lcd_nrst_s1_begins_xfer;
  wire             tft_lcd_nrst_s1_chipselect;
  wire    [  3: 0] tft_lcd_nrst_s1_chosen_master_double_vector;
  wire    [  1: 0] tft_lcd_nrst_s1_chosen_master_rot_left;
  wire             tft_lcd_nrst_s1_end_xfer;
  wire             tft_lcd_nrst_s1_firsttransfer;
  wire    [  1: 0] tft_lcd_nrst_s1_grant_vector;
  wire             tft_lcd_nrst_s1_in_a_read_cycle;
  wire             tft_lcd_nrst_s1_in_a_write_cycle;
  wire    [  1: 0] tft_lcd_nrst_s1_master_qreq_vector;
  wire             tft_lcd_nrst_s1_non_bursting_master_requests;
  wire             tft_lcd_nrst_s1_readdata_from_sa;
  reg              tft_lcd_nrst_s1_reg_firsttransfer;
  wire             tft_lcd_nrst_s1_reset_n;
  reg     [  1: 0] tft_lcd_nrst_s1_saved_chosen_master_vector;
  reg              tft_lcd_nrst_s1_slavearbiterlockenable;
  wire             tft_lcd_nrst_s1_slavearbiterlockenable2;
  wire             tft_lcd_nrst_s1_unreg_firsttransfer;
  wire             tft_lcd_nrst_s1_waits_for_read;
  wire             tft_lcd_nrst_s1_waits_for_write;
  wire             tft_lcd_nrst_s1_write_n;
  wire             tft_lcd_nrst_s1_writedata;
  wire             wait_for_tft_lcd_nrst_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tft_lcd_nrst_s1_end_xfer;
    end


  assign tft_lcd_nrst_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 | cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1));
  //assign tft_lcd_nrst_s1_readdata_from_sa = tft_lcd_nrst_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tft_lcd_nrst_s1_readdata_from_sa = tft_lcd_nrst_s1_readdata;

  assign cpu_0_data_master_requests_tft_lcd_nrst_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801080) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //tft_lcd_nrst_s1_arb_share_counter set values, which is an e_mux
  assign tft_lcd_nrst_s1_arb_share_set_values = 1;

  //tft_lcd_nrst_s1_non_bursting_master_requests mux, which is an e_mux
  assign tft_lcd_nrst_s1_non_bursting_master_requests = cpu_0_data_master_requests_tft_lcd_nrst_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nrst_s1 |
    cpu_0_data_master_requests_tft_lcd_nrst_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nrst_s1;

  //tft_lcd_nrst_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tft_lcd_nrst_s1_any_bursting_master_saved_grant = 0;

  //tft_lcd_nrst_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tft_lcd_nrst_s1_arb_share_counter_next_value = tft_lcd_nrst_s1_firsttransfer ? (tft_lcd_nrst_s1_arb_share_set_values - 1) : |tft_lcd_nrst_s1_arb_share_counter ? (tft_lcd_nrst_s1_arb_share_counter - 1) : 0;

  //tft_lcd_nrst_s1_allgrants all slave grants, which is an e_mux
  assign tft_lcd_nrst_s1_allgrants = (|tft_lcd_nrst_s1_grant_vector) |
    (|tft_lcd_nrst_s1_grant_vector) |
    (|tft_lcd_nrst_s1_grant_vector) |
    (|tft_lcd_nrst_s1_grant_vector);

  //tft_lcd_nrst_s1_end_xfer assignment, which is an e_assign
  assign tft_lcd_nrst_s1_end_xfer = ~(tft_lcd_nrst_s1_waits_for_read | tft_lcd_nrst_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tft_lcd_nrst_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tft_lcd_nrst_s1 = tft_lcd_nrst_s1_end_xfer & (~tft_lcd_nrst_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tft_lcd_nrst_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tft_lcd_nrst_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tft_lcd_nrst_s1 & tft_lcd_nrst_s1_allgrants) | (end_xfer_arb_share_counter_term_tft_lcd_nrst_s1 & ~tft_lcd_nrst_s1_non_bursting_master_requests);

  //tft_lcd_nrst_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrst_s1_arb_share_counter <= 0;
      else if (tft_lcd_nrst_s1_arb_counter_enable)
          tft_lcd_nrst_s1_arb_share_counter <= tft_lcd_nrst_s1_arb_share_counter_next_value;
    end


  //tft_lcd_nrst_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrst_s1_slavearbiterlockenable <= 0;
      else if ((|tft_lcd_nrst_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tft_lcd_nrst_s1) | (end_xfer_arb_share_counter_term_tft_lcd_nrst_s1 & ~tft_lcd_nrst_s1_non_bursting_master_requests))
          tft_lcd_nrst_s1_slavearbiterlockenable <= |tft_lcd_nrst_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master tft_lcd_nrst/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tft_lcd_nrst_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tft_lcd_nrst_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tft_lcd_nrst_s1_slavearbiterlockenable2 = |tft_lcd_nrst_s1_arb_share_counter_next_value;

  //cpu_0/data_master tft_lcd_nrst/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tft_lcd_nrst_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nrst/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tft_lcd_nrst_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nrst/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tft_lcd_nrst_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted tft_lcd_nrst/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrst_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrst_s1 <= cpu_0_instruction_master_saved_grant_tft_lcd_nrst_s1 ? 1 : (tft_lcd_nrst_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_tft_lcd_nrst_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrst_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nrst_s1 & cpu_0_instruction_master_requests_tft_lcd_nrst_s1;

  //tft_lcd_nrst_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tft_lcd_nrst_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_tft_lcd_nrst_s1 = cpu_0_data_master_requests_tft_lcd_nrst_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1 = cpu_0_data_master_granted_tft_lcd_nrst_s1 & cpu_0_data_master_read & ~tft_lcd_nrst_s1_waits_for_read;

  //tft_lcd_nrst_s1_writedata mux, which is an e_mux
  assign tft_lcd_nrst_s1_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_tft_lcd_nrst_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801080) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted tft_lcd_nrst/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrst_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrst_s1 <= cpu_0_data_master_saved_grant_tft_lcd_nrst_s1 ? 1 : (tft_lcd_nrst_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_tft_lcd_nrst_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrst_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nrst_s1 & cpu_0_data_master_requests_tft_lcd_nrst_s1;

  assign cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1 = cpu_0_instruction_master_requests_tft_lcd_nrst_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1 = cpu_0_instruction_master_granted_tft_lcd_nrst_s1 & cpu_0_instruction_master_read & ~tft_lcd_nrst_s1_waits_for_read;

  //allow new arb cycle for tft_lcd_nrst/s1, which is an e_assign
  assign tft_lcd_nrst_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for tft_lcd_nrst/s1, which is an e_assign
  assign tft_lcd_nrst_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1;

  //cpu_0/instruction_master grant tft_lcd_nrst/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_tft_lcd_nrst_s1 = tft_lcd_nrst_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant tft_lcd_nrst/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_tft_lcd_nrst_s1 = tft_lcd_nrst_s1_arb_winner[0] && cpu_0_instruction_master_requests_tft_lcd_nrst_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for tft_lcd_nrst/s1, which is an e_assign
  assign tft_lcd_nrst_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_tft_lcd_nrst_s1;

  //cpu_0/data_master grant tft_lcd_nrst/s1, which is an e_assign
  assign cpu_0_data_master_granted_tft_lcd_nrst_s1 = tft_lcd_nrst_s1_grant_vector[1];

  //cpu_0/data_master saved-grant tft_lcd_nrst/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_tft_lcd_nrst_s1 = tft_lcd_nrst_s1_arb_winner[1] && cpu_0_data_master_requests_tft_lcd_nrst_s1;

  //tft_lcd_nrst/s1 chosen-master double-vector, which is an e_assign
  assign tft_lcd_nrst_s1_chosen_master_double_vector = {tft_lcd_nrst_s1_master_qreq_vector, tft_lcd_nrst_s1_master_qreq_vector} & ({~tft_lcd_nrst_s1_master_qreq_vector, ~tft_lcd_nrst_s1_master_qreq_vector} + tft_lcd_nrst_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign tft_lcd_nrst_s1_arb_winner = (tft_lcd_nrst_s1_allow_new_arb_cycle & | tft_lcd_nrst_s1_grant_vector) ? tft_lcd_nrst_s1_grant_vector : tft_lcd_nrst_s1_saved_chosen_master_vector;

  //saved tft_lcd_nrst_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrst_s1_saved_chosen_master_vector <= 0;
      else if (tft_lcd_nrst_s1_allow_new_arb_cycle)
          tft_lcd_nrst_s1_saved_chosen_master_vector <= |tft_lcd_nrst_s1_grant_vector ? tft_lcd_nrst_s1_grant_vector : tft_lcd_nrst_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tft_lcd_nrst_s1_grant_vector = {(tft_lcd_nrst_s1_chosen_master_double_vector[1] | tft_lcd_nrst_s1_chosen_master_double_vector[3]),
    (tft_lcd_nrst_s1_chosen_master_double_vector[0] | tft_lcd_nrst_s1_chosen_master_double_vector[2])};

  //tft_lcd_nrst/s1 chosen master rotated left, which is an e_assign
  assign tft_lcd_nrst_s1_chosen_master_rot_left = (tft_lcd_nrst_s1_arb_winner << 1) ? (tft_lcd_nrst_s1_arb_winner << 1) : 1;

  //tft_lcd_nrst/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrst_s1_arb_addend <= 1;
      else if (|tft_lcd_nrst_s1_grant_vector)
          tft_lcd_nrst_s1_arb_addend <= tft_lcd_nrst_s1_end_xfer? tft_lcd_nrst_s1_chosen_master_rot_left : tft_lcd_nrst_s1_grant_vector;
    end


  //tft_lcd_nrst_s1_reset_n assignment, which is an e_assign
  assign tft_lcd_nrst_s1_reset_n = reset_n;

  assign tft_lcd_nrst_s1_chipselect = cpu_0_data_master_granted_tft_lcd_nrst_s1 | cpu_0_instruction_master_granted_tft_lcd_nrst_s1;
  //tft_lcd_nrst_s1_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nrst_s1_firsttransfer = tft_lcd_nrst_s1_begins_xfer ? tft_lcd_nrst_s1_unreg_firsttransfer : tft_lcd_nrst_s1_reg_firsttransfer;

  //tft_lcd_nrst_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nrst_s1_unreg_firsttransfer = ~(tft_lcd_nrst_s1_slavearbiterlockenable & tft_lcd_nrst_s1_any_continuerequest);

  //tft_lcd_nrst_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nrst_s1_reg_firsttransfer <= 1'b1;
      else if (tft_lcd_nrst_s1_begins_xfer)
          tft_lcd_nrst_s1_reg_firsttransfer <= tft_lcd_nrst_s1_unreg_firsttransfer;
    end


  //tft_lcd_nrst_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tft_lcd_nrst_s1_beginbursttransfer_internal = tft_lcd_nrst_s1_begins_xfer;

  //tft_lcd_nrst_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tft_lcd_nrst_s1_arbitration_holdoff_internal = tft_lcd_nrst_s1_begins_xfer & tft_lcd_nrst_s1_firsttransfer;

  //~tft_lcd_nrst_s1_write_n assignment, which is an e_mux
  assign tft_lcd_nrst_s1_write_n = ~(cpu_0_data_master_granted_tft_lcd_nrst_s1 & cpu_0_data_master_write);

  assign shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //tft_lcd_nrst_s1_address mux, which is an e_mux
  assign tft_lcd_nrst_s1_address = (cpu_0_data_master_granted_tft_lcd_nrst_s1)? (shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_data_master >> 2) :
    (shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_tft_lcd_nrst_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_tft_lcd_nrst_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tft_lcd_nrst_s1_end_xfer <= 1;
      else 
        d1_tft_lcd_nrst_s1_end_xfer <= tft_lcd_nrst_s1_end_xfer;
    end


  //tft_lcd_nrst_s1_waits_for_read in a cycle, which is an e_mux
  assign tft_lcd_nrst_s1_waits_for_read = tft_lcd_nrst_s1_in_a_read_cycle & tft_lcd_nrst_s1_begins_xfer;

  //tft_lcd_nrst_s1_in_a_read_cycle assignment, which is an e_assign
  assign tft_lcd_nrst_s1_in_a_read_cycle = (cpu_0_data_master_granted_tft_lcd_nrst_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_tft_lcd_nrst_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tft_lcd_nrst_s1_in_a_read_cycle;

  //tft_lcd_nrst_s1_waits_for_write in a cycle, which is an e_mux
  assign tft_lcd_nrst_s1_waits_for_write = tft_lcd_nrst_s1_in_a_write_cycle & 0;

  //tft_lcd_nrst_s1_in_a_write_cycle assignment, which is an e_assign
  assign tft_lcd_nrst_s1_in_a_write_cycle = cpu_0_data_master_granted_tft_lcd_nrst_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tft_lcd_nrst_s1_in_a_write_cycle;

  assign wait_for_tft_lcd_nrst_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tft_lcd_nrst/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_tft_lcd_nrst_s1 + cpu_0_instruction_master_granted_tft_lcd_nrst_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_tft_lcd_nrst_s1 + cpu_0_instruction_master_saved_grant_tft_lcd_nrst_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tft_lcd_nwr_s1_arbitrator (
                                   // inputs:
                                    clk,
                                    cpu_0_data_master_address_to_slave,
                                    cpu_0_data_master_latency_counter,
                                    cpu_0_data_master_read,
                                    cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                    cpu_0_data_master_write,
                                    cpu_0_data_master_writedata,
                                    cpu_0_instruction_master_address_to_slave,
                                    cpu_0_instruction_master_latency_counter,
                                    cpu_0_instruction_master_read,
                                    cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                    reset_n,
                                    tft_lcd_nwr_s1_readdata,

                                   // outputs:
                                    cpu_0_data_master_granted_tft_lcd_nwr_s1,
                                    cpu_0_data_master_qualified_request_tft_lcd_nwr_s1,
                                    cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1,
                                    cpu_0_data_master_requests_tft_lcd_nwr_s1,
                                    cpu_0_instruction_master_granted_tft_lcd_nwr_s1,
                                    cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1,
                                    cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1,
                                    cpu_0_instruction_master_requests_tft_lcd_nwr_s1,
                                    d1_tft_lcd_nwr_s1_end_xfer,
                                    tft_lcd_nwr_s1_address,
                                    tft_lcd_nwr_s1_chipselect,
                                    tft_lcd_nwr_s1_readdata_from_sa,
                                    tft_lcd_nwr_s1_reset_n,
                                    tft_lcd_nwr_s1_write_n,
                                    tft_lcd_nwr_s1_writedata
                                 )
;

  output           cpu_0_data_master_granted_tft_lcd_nwr_s1;
  output           cpu_0_data_master_qualified_request_tft_lcd_nwr_s1;
  output           cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1;
  output           cpu_0_data_master_requests_tft_lcd_nwr_s1;
  output           cpu_0_instruction_master_granted_tft_lcd_nwr_s1;
  output           cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1;
  output           cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1;
  output           cpu_0_instruction_master_requests_tft_lcd_nwr_s1;
  output           d1_tft_lcd_nwr_s1_end_xfer;
  output  [  1: 0] tft_lcd_nwr_s1_address;
  output           tft_lcd_nwr_s1_chipselect;
  output           tft_lcd_nwr_s1_readdata_from_sa;
  output           tft_lcd_nwr_s1_reset_n;
  output           tft_lcd_nwr_s1_write_n;
  output           tft_lcd_nwr_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;
  input            tft_lcd_nwr_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_saved_grant_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_saved_grant_tft_lcd_nwr_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tft_lcd_nwr_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tft_lcd_nwr_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nwr_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nwr_s1;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_instruction_master;
  wire    [  1: 0] tft_lcd_nwr_s1_address;
  wire             tft_lcd_nwr_s1_allgrants;
  wire             tft_lcd_nwr_s1_allow_new_arb_cycle;
  wire             tft_lcd_nwr_s1_any_bursting_master_saved_grant;
  wire             tft_lcd_nwr_s1_any_continuerequest;
  reg     [  1: 0] tft_lcd_nwr_s1_arb_addend;
  wire             tft_lcd_nwr_s1_arb_counter_enable;
  reg     [  1: 0] tft_lcd_nwr_s1_arb_share_counter;
  wire    [  1: 0] tft_lcd_nwr_s1_arb_share_counter_next_value;
  wire    [  1: 0] tft_lcd_nwr_s1_arb_share_set_values;
  wire    [  1: 0] tft_lcd_nwr_s1_arb_winner;
  wire             tft_lcd_nwr_s1_arbitration_holdoff_internal;
  wire             tft_lcd_nwr_s1_beginbursttransfer_internal;
  wire             tft_lcd_nwr_s1_begins_xfer;
  wire             tft_lcd_nwr_s1_chipselect;
  wire    [  3: 0] tft_lcd_nwr_s1_chosen_master_double_vector;
  wire    [  1: 0] tft_lcd_nwr_s1_chosen_master_rot_left;
  wire             tft_lcd_nwr_s1_end_xfer;
  wire             tft_lcd_nwr_s1_firsttransfer;
  wire    [  1: 0] tft_lcd_nwr_s1_grant_vector;
  wire             tft_lcd_nwr_s1_in_a_read_cycle;
  wire             tft_lcd_nwr_s1_in_a_write_cycle;
  wire    [  1: 0] tft_lcd_nwr_s1_master_qreq_vector;
  wire             tft_lcd_nwr_s1_non_bursting_master_requests;
  wire             tft_lcd_nwr_s1_readdata_from_sa;
  reg              tft_lcd_nwr_s1_reg_firsttransfer;
  wire             tft_lcd_nwr_s1_reset_n;
  reg     [  1: 0] tft_lcd_nwr_s1_saved_chosen_master_vector;
  reg              tft_lcd_nwr_s1_slavearbiterlockenable;
  wire             tft_lcd_nwr_s1_slavearbiterlockenable2;
  wire             tft_lcd_nwr_s1_unreg_firsttransfer;
  wire             tft_lcd_nwr_s1_waits_for_read;
  wire             tft_lcd_nwr_s1_waits_for_write;
  wire             tft_lcd_nwr_s1_write_n;
  wire             tft_lcd_nwr_s1_writedata;
  wire             wait_for_tft_lcd_nwr_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tft_lcd_nwr_s1_end_xfer;
    end


  assign tft_lcd_nwr_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 | cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1));
  //assign tft_lcd_nwr_s1_readdata_from_sa = tft_lcd_nwr_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tft_lcd_nwr_s1_readdata_from_sa = tft_lcd_nwr_s1_readdata;

  assign cpu_0_data_master_requests_tft_lcd_nwr_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010b0) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //tft_lcd_nwr_s1_arb_share_counter set values, which is an e_mux
  assign tft_lcd_nwr_s1_arb_share_set_values = 1;

  //tft_lcd_nwr_s1_non_bursting_master_requests mux, which is an e_mux
  assign tft_lcd_nwr_s1_non_bursting_master_requests = cpu_0_data_master_requests_tft_lcd_nwr_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nwr_s1 |
    cpu_0_data_master_requests_tft_lcd_nwr_s1 |
    cpu_0_instruction_master_requests_tft_lcd_nwr_s1;

  //tft_lcd_nwr_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tft_lcd_nwr_s1_any_bursting_master_saved_grant = 0;

  //tft_lcd_nwr_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tft_lcd_nwr_s1_arb_share_counter_next_value = tft_lcd_nwr_s1_firsttransfer ? (tft_lcd_nwr_s1_arb_share_set_values - 1) : |tft_lcd_nwr_s1_arb_share_counter ? (tft_lcd_nwr_s1_arb_share_counter - 1) : 0;

  //tft_lcd_nwr_s1_allgrants all slave grants, which is an e_mux
  assign tft_lcd_nwr_s1_allgrants = (|tft_lcd_nwr_s1_grant_vector) |
    (|tft_lcd_nwr_s1_grant_vector) |
    (|tft_lcd_nwr_s1_grant_vector) |
    (|tft_lcd_nwr_s1_grant_vector);

  //tft_lcd_nwr_s1_end_xfer assignment, which is an e_assign
  assign tft_lcd_nwr_s1_end_xfer = ~(tft_lcd_nwr_s1_waits_for_read | tft_lcd_nwr_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tft_lcd_nwr_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tft_lcd_nwr_s1 = tft_lcd_nwr_s1_end_xfer & (~tft_lcd_nwr_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tft_lcd_nwr_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tft_lcd_nwr_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tft_lcd_nwr_s1 & tft_lcd_nwr_s1_allgrants) | (end_xfer_arb_share_counter_term_tft_lcd_nwr_s1 & ~tft_lcd_nwr_s1_non_bursting_master_requests);

  //tft_lcd_nwr_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nwr_s1_arb_share_counter <= 0;
      else if (tft_lcd_nwr_s1_arb_counter_enable)
          tft_lcd_nwr_s1_arb_share_counter <= tft_lcd_nwr_s1_arb_share_counter_next_value;
    end


  //tft_lcd_nwr_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nwr_s1_slavearbiterlockenable <= 0;
      else if ((|tft_lcd_nwr_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tft_lcd_nwr_s1) | (end_xfer_arb_share_counter_term_tft_lcd_nwr_s1 & ~tft_lcd_nwr_s1_non_bursting_master_requests))
          tft_lcd_nwr_s1_slavearbiterlockenable <= |tft_lcd_nwr_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master tft_lcd_nwr/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tft_lcd_nwr_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tft_lcd_nwr_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tft_lcd_nwr_s1_slavearbiterlockenable2 = |tft_lcd_nwr_s1_arb_share_counter_next_value;

  //cpu_0/data_master tft_lcd_nwr/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tft_lcd_nwr_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nwr/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tft_lcd_nwr_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_nwr/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tft_lcd_nwr_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted tft_lcd_nwr/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nwr_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nwr_s1 <= cpu_0_instruction_master_saved_grant_tft_lcd_nwr_s1 ? 1 : (tft_lcd_nwr_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_tft_lcd_nwr_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nwr_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_nwr_s1 & cpu_0_instruction_master_requests_tft_lcd_nwr_s1;

  //tft_lcd_nwr_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tft_lcd_nwr_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_tft_lcd_nwr_s1 = cpu_0_data_master_requests_tft_lcd_nwr_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1 = cpu_0_data_master_granted_tft_lcd_nwr_s1 & cpu_0_data_master_read & ~tft_lcd_nwr_s1_waits_for_read;

  //tft_lcd_nwr_s1_writedata mux, which is an e_mux
  assign tft_lcd_nwr_s1_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_tft_lcd_nwr_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 4] , 4'b0} == 25'h18010b0) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted tft_lcd_nwr/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nwr_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nwr_s1 <= cpu_0_data_master_saved_grant_tft_lcd_nwr_s1 ? 1 : (tft_lcd_nwr_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_tft_lcd_nwr_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nwr_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_tft_lcd_nwr_s1 & cpu_0_data_master_requests_tft_lcd_nwr_s1;

  assign cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1 = cpu_0_instruction_master_requests_tft_lcd_nwr_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1 = cpu_0_instruction_master_granted_tft_lcd_nwr_s1 & cpu_0_instruction_master_read & ~tft_lcd_nwr_s1_waits_for_read;

  //allow new arb cycle for tft_lcd_nwr/s1, which is an e_assign
  assign tft_lcd_nwr_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for tft_lcd_nwr/s1, which is an e_assign
  assign tft_lcd_nwr_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1;

  //cpu_0/instruction_master grant tft_lcd_nwr/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_tft_lcd_nwr_s1 = tft_lcd_nwr_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant tft_lcd_nwr/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_tft_lcd_nwr_s1 = tft_lcd_nwr_s1_arb_winner[0] && cpu_0_instruction_master_requests_tft_lcd_nwr_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for tft_lcd_nwr/s1, which is an e_assign
  assign tft_lcd_nwr_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_tft_lcd_nwr_s1;

  //cpu_0/data_master grant tft_lcd_nwr/s1, which is an e_assign
  assign cpu_0_data_master_granted_tft_lcd_nwr_s1 = tft_lcd_nwr_s1_grant_vector[1];

  //cpu_0/data_master saved-grant tft_lcd_nwr/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_tft_lcd_nwr_s1 = tft_lcd_nwr_s1_arb_winner[1] && cpu_0_data_master_requests_tft_lcd_nwr_s1;

  //tft_lcd_nwr/s1 chosen-master double-vector, which is an e_assign
  assign tft_lcd_nwr_s1_chosen_master_double_vector = {tft_lcd_nwr_s1_master_qreq_vector, tft_lcd_nwr_s1_master_qreq_vector} & ({~tft_lcd_nwr_s1_master_qreq_vector, ~tft_lcd_nwr_s1_master_qreq_vector} + tft_lcd_nwr_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign tft_lcd_nwr_s1_arb_winner = (tft_lcd_nwr_s1_allow_new_arb_cycle & | tft_lcd_nwr_s1_grant_vector) ? tft_lcd_nwr_s1_grant_vector : tft_lcd_nwr_s1_saved_chosen_master_vector;

  //saved tft_lcd_nwr_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nwr_s1_saved_chosen_master_vector <= 0;
      else if (tft_lcd_nwr_s1_allow_new_arb_cycle)
          tft_lcd_nwr_s1_saved_chosen_master_vector <= |tft_lcd_nwr_s1_grant_vector ? tft_lcd_nwr_s1_grant_vector : tft_lcd_nwr_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tft_lcd_nwr_s1_grant_vector = {(tft_lcd_nwr_s1_chosen_master_double_vector[1] | tft_lcd_nwr_s1_chosen_master_double_vector[3]),
    (tft_lcd_nwr_s1_chosen_master_double_vector[0] | tft_lcd_nwr_s1_chosen_master_double_vector[2])};

  //tft_lcd_nwr/s1 chosen master rotated left, which is an e_assign
  assign tft_lcd_nwr_s1_chosen_master_rot_left = (tft_lcd_nwr_s1_arb_winner << 1) ? (tft_lcd_nwr_s1_arb_winner << 1) : 1;

  //tft_lcd_nwr/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nwr_s1_arb_addend <= 1;
      else if (|tft_lcd_nwr_s1_grant_vector)
          tft_lcd_nwr_s1_arb_addend <= tft_lcd_nwr_s1_end_xfer? tft_lcd_nwr_s1_chosen_master_rot_left : tft_lcd_nwr_s1_grant_vector;
    end


  //tft_lcd_nwr_s1_reset_n assignment, which is an e_assign
  assign tft_lcd_nwr_s1_reset_n = reset_n;

  assign tft_lcd_nwr_s1_chipselect = cpu_0_data_master_granted_tft_lcd_nwr_s1 | cpu_0_instruction_master_granted_tft_lcd_nwr_s1;
  //tft_lcd_nwr_s1_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nwr_s1_firsttransfer = tft_lcd_nwr_s1_begins_xfer ? tft_lcd_nwr_s1_unreg_firsttransfer : tft_lcd_nwr_s1_reg_firsttransfer;

  //tft_lcd_nwr_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_nwr_s1_unreg_firsttransfer = ~(tft_lcd_nwr_s1_slavearbiterlockenable & tft_lcd_nwr_s1_any_continuerequest);

  //tft_lcd_nwr_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_nwr_s1_reg_firsttransfer <= 1'b1;
      else if (tft_lcd_nwr_s1_begins_xfer)
          tft_lcd_nwr_s1_reg_firsttransfer <= tft_lcd_nwr_s1_unreg_firsttransfer;
    end


  //tft_lcd_nwr_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tft_lcd_nwr_s1_beginbursttransfer_internal = tft_lcd_nwr_s1_begins_xfer;

  //tft_lcd_nwr_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tft_lcd_nwr_s1_arbitration_holdoff_internal = tft_lcd_nwr_s1_begins_xfer & tft_lcd_nwr_s1_firsttransfer;

  //~tft_lcd_nwr_s1_write_n assignment, which is an e_mux
  assign tft_lcd_nwr_s1_write_n = ~(cpu_0_data_master_granted_tft_lcd_nwr_s1 & cpu_0_data_master_write);

  assign shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //tft_lcd_nwr_s1_address mux, which is an e_mux
  assign tft_lcd_nwr_s1_address = (cpu_0_data_master_granted_tft_lcd_nwr_s1)? (shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_data_master >> 2) :
    (shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_tft_lcd_nwr_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_tft_lcd_nwr_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tft_lcd_nwr_s1_end_xfer <= 1;
      else 
        d1_tft_lcd_nwr_s1_end_xfer <= tft_lcd_nwr_s1_end_xfer;
    end


  //tft_lcd_nwr_s1_waits_for_read in a cycle, which is an e_mux
  assign tft_lcd_nwr_s1_waits_for_read = tft_lcd_nwr_s1_in_a_read_cycle & tft_lcd_nwr_s1_begins_xfer;

  //tft_lcd_nwr_s1_in_a_read_cycle assignment, which is an e_assign
  assign tft_lcd_nwr_s1_in_a_read_cycle = (cpu_0_data_master_granted_tft_lcd_nwr_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_tft_lcd_nwr_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tft_lcd_nwr_s1_in_a_read_cycle;

  //tft_lcd_nwr_s1_waits_for_write in a cycle, which is an e_mux
  assign tft_lcd_nwr_s1_waits_for_write = tft_lcd_nwr_s1_in_a_write_cycle & 0;

  //tft_lcd_nwr_s1_in_a_write_cycle assignment, which is an e_assign
  assign tft_lcd_nwr_s1_in_a_write_cycle = cpu_0_data_master_granted_tft_lcd_nwr_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tft_lcd_nwr_s1_in_a_write_cycle;

  assign wait_for_tft_lcd_nwr_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tft_lcd_nwr/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_tft_lcd_nwr_s1 + cpu_0_instruction_master_granted_tft_lcd_nwr_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_tft_lcd_nwr_s1 + cpu_0_instruction_master_saved_grant_tft_lcd_nwr_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tft_lcd_rs_s1_arbitrator (
                                  // inputs:
                                   clk,
                                   cpu_0_data_master_address_to_slave,
                                   cpu_0_data_master_latency_counter,
                                   cpu_0_data_master_read,
                                   cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                   cpu_0_data_master_write,
                                   cpu_0_data_master_writedata,
                                   cpu_0_instruction_master_address_to_slave,
                                   cpu_0_instruction_master_latency_counter,
                                   cpu_0_instruction_master_read,
                                   cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                   reset_n,
                                   tft_lcd_rs_s1_readdata,

                                  // outputs:
                                   cpu_0_data_master_granted_tft_lcd_rs_s1,
                                   cpu_0_data_master_qualified_request_tft_lcd_rs_s1,
                                   cpu_0_data_master_read_data_valid_tft_lcd_rs_s1,
                                   cpu_0_data_master_requests_tft_lcd_rs_s1,
                                   cpu_0_instruction_master_granted_tft_lcd_rs_s1,
                                   cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1,
                                   cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1,
                                   cpu_0_instruction_master_requests_tft_lcd_rs_s1,
                                   d1_tft_lcd_rs_s1_end_xfer,
                                   tft_lcd_rs_s1_address,
                                   tft_lcd_rs_s1_chipselect,
                                   tft_lcd_rs_s1_readdata_from_sa,
                                   tft_lcd_rs_s1_reset_n,
                                   tft_lcd_rs_s1_write_n,
                                   tft_lcd_rs_s1_writedata
                                )
;

  output           cpu_0_data_master_granted_tft_lcd_rs_s1;
  output           cpu_0_data_master_qualified_request_tft_lcd_rs_s1;
  output           cpu_0_data_master_read_data_valid_tft_lcd_rs_s1;
  output           cpu_0_data_master_requests_tft_lcd_rs_s1;
  output           cpu_0_instruction_master_granted_tft_lcd_rs_s1;
  output           cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1;
  output           cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1;
  output           cpu_0_instruction_master_requests_tft_lcd_rs_s1;
  output           d1_tft_lcd_rs_s1_end_xfer;
  output  [  1: 0] tft_lcd_rs_s1_address;
  output           tft_lcd_rs_s1_chipselect;
  output           tft_lcd_rs_s1_readdata_from_sa;
  output           tft_lcd_rs_s1_reset_n;
  output           tft_lcd_rs_s1_write_n;
  output           tft_lcd_rs_s1_writedata;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 31: 0] cpu_0_data_master_writedata;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;
  input            tft_lcd_rs_s1_readdata;

  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_tft_lcd_rs_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_rs_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_rs_s1;
  wire             cpu_0_data_master_requests_tft_lcd_rs_s1;
  wire             cpu_0_data_master_saved_grant_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_saved_grant_tft_lcd_rs_s1;
  reg              d1_reasons_to_wait;
  reg              d1_tft_lcd_rs_s1_end_xfer;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tft_lcd_rs_s1;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg              last_cycle_cpu_0_data_master_granted_slave_tft_lcd_rs_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_rs_s1;
  wire    [ 24: 0] shifted_address_to_tft_lcd_rs_s1_from_cpu_0_data_master;
  wire    [ 24: 0] shifted_address_to_tft_lcd_rs_s1_from_cpu_0_instruction_master;
  wire    [  1: 0] tft_lcd_rs_s1_address;
  wire             tft_lcd_rs_s1_allgrants;
  wire             tft_lcd_rs_s1_allow_new_arb_cycle;
  wire             tft_lcd_rs_s1_any_bursting_master_saved_grant;
  wire             tft_lcd_rs_s1_any_continuerequest;
  reg     [  1: 0] tft_lcd_rs_s1_arb_addend;
  wire             tft_lcd_rs_s1_arb_counter_enable;
  reg     [  1: 0] tft_lcd_rs_s1_arb_share_counter;
  wire    [  1: 0] tft_lcd_rs_s1_arb_share_counter_next_value;
  wire    [  1: 0] tft_lcd_rs_s1_arb_share_set_values;
  wire    [  1: 0] tft_lcd_rs_s1_arb_winner;
  wire             tft_lcd_rs_s1_arbitration_holdoff_internal;
  wire             tft_lcd_rs_s1_beginbursttransfer_internal;
  wire             tft_lcd_rs_s1_begins_xfer;
  wire             tft_lcd_rs_s1_chipselect;
  wire    [  3: 0] tft_lcd_rs_s1_chosen_master_double_vector;
  wire    [  1: 0] tft_lcd_rs_s1_chosen_master_rot_left;
  wire             tft_lcd_rs_s1_end_xfer;
  wire             tft_lcd_rs_s1_firsttransfer;
  wire    [  1: 0] tft_lcd_rs_s1_grant_vector;
  wire             tft_lcd_rs_s1_in_a_read_cycle;
  wire             tft_lcd_rs_s1_in_a_write_cycle;
  wire    [  1: 0] tft_lcd_rs_s1_master_qreq_vector;
  wire             tft_lcd_rs_s1_non_bursting_master_requests;
  wire             tft_lcd_rs_s1_readdata_from_sa;
  reg              tft_lcd_rs_s1_reg_firsttransfer;
  wire             tft_lcd_rs_s1_reset_n;
  reg     [  1: 0] tft_lcd_rs_s1_saved_chosen_master_vector;
  reg              tft_lcd_rs_s1_slavearbiterlockenable;
  wire             tft_lcd_rs_s1_slavearbiterlockenable2;
  wire             tft_lcd_rs_s1_unreg_firsttransfer;
  wire             tft_lcd_rs_s1_waits_for_read;
  wire             tft_lcd_rs_s1_waits_for_write;
  wire             tft_lcd_rs_s1_write_n;
  wire             tft_lcd_rs_s1_writedata;
  wire             wait_for_tft_lcd_rs_s1_counter;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tft_lcd_rs_s1_end_xfer;
    end


  assign tft_lcd_rs_s1_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_tft_lcd_rs_s1 | cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1));
  //assign tft_lcd_rs_s1_readdata_from_sa = tft_lcd_rs_s1_readdata so that symbol knows where to group signals which may go to master only, which is an e_assign
  assign tft_lcd_rs_s1_readdata_from_sa = tft_lcd_rs_s1_readdata;

  assign cpu_0_data_master_requests_tft_lcd_rs_s1 = ({cpu_0_data_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801090) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //tft_lcd_rs_s1_arb_share_counter set values, which is an e_mux
  assign tft_lcd_rs_s1_arb_share_set_values = 1;

  //tft_lcd_rs_s1_non_bursting_master_requests mux, which is an e_mux
  assign tft_lcd_rs_s1_non_bursting_master_requests = cpu_0_data_master_requests_tft_lcd_rs_s1 |
    cpu_0_instruction_master_requests_tft_lcd_rs_s1 |
    cpu_0_data_master_requests_tft_lcd_rs_s1 |
    cpu_0_instruction_master_requests_tft_lcd_rs_s1;

  //tft_lcd_rs_s1_any_bursting_master_saved_grant mux, which is an e_mux
  assign tft_lcd_rs_s1_any_bursting_master_saved_grant = 0;

  //tft_lcd_rs_s1_arb_share_counter_next_value assignment, which is an e_assign
  assign tft_lcd_rs_s1_arb_share_counter_next_value = tft_lcd_rs_s1_firsttransfer ? (tft_lcd_rs_s1_arb_share_set_values - 1) : |tft_lcd_rs_s1_arb_share_counter ? (tft_lcd_rs_s1_arb_share_counter - 1) : 0;

  //tft_lcd_rs_s1_allgrants all slave grants, which is an e_mux
  assign tft_lcd_rs_s1_allgrants = (|tft_lcd_rs_s1_grant_vector) |
    (|tft_lcd_rs_s1_grant_vector) |
    (|tft_lcd_rs_s1_grant_vector) |
    (|tft_lcd_rs_s1_grant_vector);

  //tft_lcd_rs_s1_end_xfer assignment, which is an e_assign
  assign tft_lcd_rs_s1_end_xfer = ~(tft_lcd_rs_s1_waits_for_read | tft_lcd_rs_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tft_lcd_rs_s1 arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tft_lcd_rs_s1 = tft_lcd_rs_s1_end_xfer & (~tft_lcd_rs_s1_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tft_lcd_rs_s1_arb_share_counter arbitration counter enable, which is an e_assign
  assign tft_lcd_rs_s1_arb_counter_enable = (end_xfer_arb_share_counter_term_tft_lcd_rs_s1 & tft_lcd_rs_s1_allgrants) | (end_xfer_arb_share_counter_term_tft_lcd_rs_s1 & ~tft_lcd_rs_s1_non_bursting_master_requests);

  //tft_lcd_rs_s1_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_rs_s1_arb_share_counter <= 0;
      else if (tft_lcd_rs_s1_arb_counter_enable)
          tft_lcd_rs_s1_arb_share_counter <= tft_lcd_rs_s1_arb_share_counter_next_value;
    end


  //tft_lcd_rs_s1_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_rs_s1_slavearbiterlockenable <= 0;
      else if ((|tft_lcd_rs_s1_master_qreq_vector & end_xfer_arb_share_counter_term_tft_lcd_rs_s1) | (end_xfer_arb_share_counter_term_tft_lcd_rs_s1 & ~tft_lcd_rs_s1_non_bursting_master_requests))
          tft_lcd_rs_s1_slavearbiterlockenable <= |tft_lcd_rs_s1_arb_share_counter_next_value;
    end


  //cpu_0/data_master tft_lcd_rs/s1 arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tft_lcd_rs_s1_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tft_lcd_rs_s1_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tft_lcd_rs_s1_slavearbiterlockenable2 = |tft_lcd_rs_s1_arb_share_counter_next_value;

  //cpu_0/data_master tft_lcd_rs/s1 arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tft_lcd_rs_s1_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_rs/s1 arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tft_lcd_rs_s1_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tft_lcd_rs/s1 arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tft_lcd_rs_s1_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted tft_lcd_rs/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_rs_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_rs_s1 <= cpu_0_instruction_master_saved_grant_tft_lcd_rs_s1 ? 1 : (tft_lcd_rs_s1_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_tft_lcd_rs_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_rs_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_tft_lcd_rs_s1 & cpu_0_instruction_master_requests_tft_lcd_rs_s1;

  //tft_lcd_rs_s1_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tft_lcd_rs_s1_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_tft_lcd_rs_s1 = cpu_0_data_master_requests_tft_lcd_rs_s1 & ~((cpu_0_data_master_read & ((cpu_0_data_master_latency_counter != 0) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_instruction_master_arbiterlock);
  //local readdatavalid cpu_0_data_master_read_data_valid_tft_lcd_rs_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_tft_lcd_rs_s1 = cpu_0_data_master_granted_tft_lcd_rs_s1 & cpu_0_data_master_read & ~tft_lcd_rs_s1_waits_for_read;

  //tft_lcd_rs_s1_writedata mux, which is an e_mux
  assign tft_lcd_rs_s1_writedata = cpu_0_data_master_writedata;

  assign cpu_0_instruction_master_requests_tft_lcd_rs_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 4] , 4'b0} == 25'h1801090) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted tft_lcd_rs/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_tft_lcd_rs_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_tft_lcd_rs_s1 <= cpu_0_data_master_saved_grant_tft_lcd_rs_s1 ? 1 : (tft_lcd_rs_s1_arbitration_holdoff_internal | ~cpu_0_data_master_requests_tft_lcd_rs_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_tft_lcd_rs_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_tft_lcd_rs_s1 & cpu_0_data_master_requests_tft_lcd_rs_s1;

  assign cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1 = cpu_0_instruction_master_requests_tft_lcd_rs_s1 & ~((cpu_0_instruction_master_read & ((cpu_0_instruction_master_latency_counter != 0) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //local readdatavalid cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1 = cpu_0_instruction_master_granted_tft_lcd_rs_s1 & cpu_0_instruction_master_read & ~tft_lcd_rs_s1_waits_for_read;

  //allow new arb cycle for tft_lcd_rs/s1, which is an e_assign
  assign tft_lcd_rs_s1_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for tft_lcd_rs/s1, which is an e_assign
  assign tft_lcd_rs_s1_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1;

  //cpu_0/instruction_master grant tft_lcd_rs/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_tft_lcd_rs_s1 = tft_lcd_rs_s1_grant_vector[0];

  //cpu_0/instruction_master saved-grant tft_lcd_rs/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_tft_lcd_rs_s1 = tft_lcd_rs_s1_arb_winner[0] && cpu_0_instruction_master_requests_tft_lcd_rs_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for tft_lcd_rs/s1, which is an e_assign
  assign tft_lcd_rs_s1_master_qreq_vector[1] = cpu_0_data_master_qualified_request_tft_lcd_rs_s1;

  //cpu_0/data_master grant tft_lcd_rs/s1, which is an e_assign
  assign cpu_0_data_master_granted_tft_lcd_rs_s1 = tft_lcd_rs_s1_grant_vector[1];

  //cpu_0/data_master saved-grant tft_lcd_rs/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_tft_lcd_rs_s1 = tft_lcd_rs_s1_arb_winner[1] && cpu_0_data_master_requests_tft_lcd_rs_s1;

  //tft_lcd_rs/s1 chosen-master double-vector, which is an e_assign
  assign tft_lcd_rs_s1_chosen_master_double_vector = {tft_lcd_rs_s1_master_qreq_vector, tft_lcd_rs_s1_master_qreq_vector} & ({~tft_lcd_rs_s1_master_qreq_vector, ~tft_lcd_rs_s1_master_qreq_vector} + tft_lcd_rs_s1_arb_addend);

  //stable onehot encoding of arb winner
  assign tft_lcd_rs_s1_arb_winner = (tft_lcd_rs_s1_allow_new_arb_cycle & | tft_lcd_rs_s1_grant_vector) ? tft_lcd_rs_s1_grant_vector : tft_lcd_rs_s1_saved_chosen_master_vector;

  //saved tft_lcd_rs_s1_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_rs_s1_saved_chosen_master_vector <= 0;
      else if (tft_lcd_rs_s1_allow_new_arb_cycle)
          tft_lcd_rs_s1_saved_chosen_master_vector <= |tft_lcd_rs_s1_grant_vector ? tft_lcd_rs_s1_grant_vector : tft_lcd_rs_s1_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tft_lcd_rs_s1_grant_vector = {(tft_lcd_rs_s1_chosen_master_double_vector[1] | tft_lcd_rs_s1_chosen_master_double_vector[3]),
    (tft_lcd_rs_s1_chosen_master_double_vector[0] | tft_lcd_rs_s1_chosen_master_double_vector[2])};

  //tft_lcd_rs/s1 chosen master rotated left, which is an e_assign
  assign tft_lcd_rs_s1_chosen_master_rot_left = (tft_lcd_rs_s1_arb_winner << 1) ? (tft_lcd_rs_s1_arb_winner << 1) : 1;

  //tft_lcd_rs/s1's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_rs_s1_arb_addend <= 1;
      else if (|tft_lcd_rs_s1_grant_vector)
          tft_lcd_rs_s1_arb_addend <= tft_lcd_rs_s1_end_xfer? tft_lcd_rs_s1_chosen_master_rot_left : tft_lcd_rs_s1_grant_vector;
    end


  //tft_lcd_rs_s1_reset_n assignment, which is an e_assign
  assign tft_lcd_rs_s1_reset_n = reset_n;

  assign tft_lcd_rs_s1_chipselect = cpu_0_data_master_granted_tft_lcd_rs_s1 | cpu_0_instruction_master_granted_tft_lcd_rs_s1;
  //tft_lcd_rs_s1_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_rs_s1_firsttransfer = tft_lcd_rs_s1_begins_xfer ? tft_lcd_rs_s1_unreg_firsttransfer : tft_lcd_rs_s1_reg_firsttransfer;

  //tft_lcd_rs_s1_unreg_firsttransfer first transaction, which is an e_assign
  assign tft_lcd_rs_s1_unreg_firsttransfer = ~(tft_lcd_rs_s1_slavearbiterlockenable & tft_lcd_rs_s1_any_continuerequest);

  //tft_lcd_rs_s1_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tft_lcd_rs_s1_reg_firsttransfer <= 1'b1;
      else if (tft_lcd_rs_s1_begins_xfer)
          tft_lcd_rs_s1_reg_firsttransfer <= tft_lcd_rs_s1_unreg_firsttransfer;
    end


  //tft_lcd_rs_s1_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tft_lcd_rs_s1_beginbursttransfer_internal = tft_lcd_rs_s1_begins_xfer;

  //tft_lcd_rs_s1_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tft_lcd_rs_s1_arbitration_holdoff_internal = tft_lcd_rs_s1_begins_xfer & tft_lcd_rs_s1_firsttransfer;

  //~tft_lcd_rs_s1_write_n assignment, which is an e_mux
  assign tft_lcd_rs_s1_write_n = ~(cpu_0_data_master_granted_tft_lcd_rs_s1 & cpu_0_data_master_write);

  assign shifted_address_to_tft_lcd_rs_s1_from_cpu_0_data_master = cpu_0_data_master_address_to_slave;
  //tft_lcd_rs_s1_address mux, which is an e_mux
  assign tft_lcd_rs_s1_address = (cpu_0_data_master_granted_tft_lcd_rs_s1)? (shifted_address_to_tft_lcd_rs_s1_from_cpu_0_data_master >> 2) :
    (shifted_address_to_tft_lcd_rs_s1_from_cpu_0_instruction_master >> 2);

  assign shifted_address_to_tft_lcd_rs_s1_from_cpu_0_instruction_master = cpu_0_instruction_master_address_to_slave;
  //d1_tft_lcd_rs_s1_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tft_lcd_rs_s1_end_xfer <= 1;
      else 
        d1_tft_lcd_rs_s1_end_xfer <= tft_lcd_rs_s1_end_xfer;
    end


  //tft_lcd_rs_s1_waits_for_read in a cycle, which is an e_mux
  assign tft_lcd_rs_s1_waits_for_read = tft_lcd_rs_s1_in_a_read_cycle & tft_lcd_rs_s1_begins_xfer;

  //tft_lcd_rs_s1_in_a_read_cycle assignment, which is an e_assign
  assign tft_lcd_rs_s1_in_a_read_cycle = (cpu_0_data_master_granted_tft_lcd_rs_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_tft_lcd_rs_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = tft_lcd_rs_s1_in_a_read_cycle;

  //tft_lcd_rs_s1_waits_for_write in a cycle, which is an e_mux
  assign tft_lcd_rs_s1_waits_for_write = tft_lcd_rs_s1_in_a_write_cycle & 0;

  //tft_lcd_rs_s1_in_a_write_cycle assignment, which is an e_assign
  assign tft_lcd_rs_s1_in_a_write_cycle = cpu_0_data_master_granted_tft_lcd_rs_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = tft_lcd_rs_s1_in_a_write_cycle;

  assign wait_for_tft_lcd_rs_s1_counter = 0;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //tft_lcd_rs/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_tft_lcd_rs_s1 + cpu_0_instruction_master_granted_tft_lcd_rs_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_tft_lcd_rs_s1 + cpu_0_instruction_master_saved_grant_tft_lcd_rs_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tri_state_bridge_0_avalon_slave_arbitrator (
                                                    // inputs:
                                                     clk,
                                                     cpu_0_data_master_address_to_slave,
                                                     cpu_0_data_master_byteenable,
                                                     cpu_0_data_master_dbs_address,
                                                     cpu_0_data_master_dbs_write_16,
                                                     cpu_0_data_master_latency_counter,
                                                     cpu_0_data_master_read,
                                                     cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register,
                                                     cpu_0_data_master_write,
                                                     cpu_0_instruction_master_address_to_slave,
                                                     cpu_0_instruction_master_dbs_address,
                                                     cpu_0_instruction_master_latency_counter,
                                                     cpu_0_instruction_master_read,
                                                     cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register,
                                                     reset_n,

                                                    // outputs:
                                                     address_to_the_cfi_flash_0,
                                                     cfi_flash_0_s1_wait_counter_eq_0,
                                                     cpu_0_data_master_byteenable_cfi_flash_0_s1,
                                                     cpu_0_data_master_granted_cfi_flash_0_s1,
                                                     cpu_0_data_master_qualified_request_cfi_flash_0_s1,
                                                     cpu_0_data_master_read_data_valid_cfi_flash_0_s1,
                                                     cpu_0_data_master_requests_cfi_flash_0_s1,
                                                     cpu_0_instruction_master_granted_cfi_flash_0_s1,
                                                     cpu_0_instruction_master_qualified_request_cfi_flash_0_s1,
                                                     cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1,
                                                     cpu_0_instruction_master_requests_cfi_flash_0_s1,
                                                     d1_tri_state_bridge_0_avalon_slave_end_xfer,
                                                     data_to_and_from_the_cfi_flash_0,
                                                     incoming_data_to_and_from_the_cfi_flash_0,
                                                     incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0,
                                                     read_n_to_the_cfi_flash_0,
                                                     select_n_to_the_cfi_flash_0,
                                                     write_n_to_the_cfi_flash_0
                                                  )
;

  output  [ 21: 0] address_to_the_cfi_flash_0;
  output           cfi_flash_0_s1_wait_counter_eq_0;
  output  [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1;
  output           cpu_0_data_master_granted_cfi_flash_0_s1;
  output           cpu_0_data_master_qualified_request_cfi_flash_0_s1;
  output           cpu_0_data_master_read_data_valid_cfi_flash_0_s1;
  output           cpu_0_data_master_requests_cfi_flash_0_s1;
  output           cpu_0_instruction_master_granted_cfi_flash_0_s1;
  output           cpu_0_instruction_master_qualified_request_cfi_flash_0_s1;
  output           cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1;
  output           cpu_0_instruction_master_requests_cfi_flash_0_s1;
  output           d1_tri_state_bridge_0_avalon_slave_end_xfer;
  inout   [ 15: 0] data_to_and_from_the_cfi_flash_0;
  output  [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0;
  output  [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0;
  output           read_n_to_the_cfi_flash_0;
  output           select_n_to_the_cfi_flash_0;
  output           write_n_to_the_cfi_flash_0;
  input            clk;
  input   [ 24: 0] cpu_0_data_master_address_to_slave;
  input   [  3: 0] cpu_0_data_master_byteenable;
  input   [  1: 0] cpu_0_data_master_dbs_address;
  input   [ 15: 0] cpu_0_data_master_dbs_write_16;
  input   [  1: 0] cpu_0_data_master_latency_counter;
  input            cpu_0_data_master_read;
  input            cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  input            cpu_0_data_master_write;
  input   [ 24: 0] cpu_0_instruction_master_address_to_slave;
  input   [  1: 0] cpu_0_instruction_master_dbs_address;
  input   [  1: 0] cpu_0_instruction_master_latency_counter;
  input            cpu_0_instruction_master_read;
  input            cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  input            reset_n;

  reg     [ 21: 0] address_to_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire    [  3: 0] cfi_flash_0_s1_counter_load_value;
  wire             cfi_flash_0_s1_in_a_read_cycle;
  wire             cfi_flash_0_s1_in_a_write_cycle;
  reg     [  3: 0] cfi_flash_0_s1_wait_counter;
  wire             cfi_flash_0_s1_wait_counter_eq_0;
  wire             cfi_flash_0_s1_waits_for_read;
  wire             cfi_flash_0_s1_waits_for_write;
  wire             cfi_flash_0_s1_with_write_latency;
  wire             cpu_0_data_master_arbiterlock;
  wire             cpu_0_data_master_arbiterlock2;
  wire    [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1;
  wire    [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_0;
  wire    [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_1;
  wire             cpu_0_data_master_continuerequest;
  wire             cpu_0_data_master_granted_cfi_flash_0_s1;
  wire             cpu_0_data_master_qualified_request_cfi_flash_0_s1;
  wire             cpu_0_data_master_read_data_valid_cfi_flash_0_s1;
  reg     [  1: 0] cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in;
  wire             cpu_0_data_master_requests_cfi_flash_0_s1;
  wire             cpu_0_data_master_saved_grant_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_arbiterlock;
  wire             cpu_0_instruction_master_arbiterlock2;
  wire             cpu_0_instruction_master_continuerequest;
  wire             cpu_0_instruction_master_granted_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_qualified_request_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1;
  reg     [  1: 0] cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in;
  wire             cpu_0_instruction_master_requests_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_saved_grant_cfi_flash_0_s1;
  reg              d1_in_a_write_cycle /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_ENABLE_REGISTER=ON"  */;
  reg     [ 15: 0] d1_outgoing_data_to_and_from_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              d1_reasons_to_wait;
  reg              d1_tri_state_bridge_0_avalon_slave_end_xfer;
  wire    [ 15: 0] data_to_and_from_the_cfi_flash_0;
  reg              enable_nonzero_assertions;
  wire             end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave;
  wire             in_a_read_cycle;
  wire             in_a_write_cycle;
  reg     [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_INPUT_REGISTER=ON"  */;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_0_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_10_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_11_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_12_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_13_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_14_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_15_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_1_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_2_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_3_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_4_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_5_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_6_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_7_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_8_is_x;
  wire             incoming_data_to_and_from_the_cfi_flash_0_bit_9_is_x;
  wire    [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0;
  reg              last_cycle_cpu_0_data_master_granted_slave_cfi_flash_0_s1;
  reg              last_cycle_cpu_0_instruction_master_granted_slave_cfi_flash_0_s1;
  wire    [ 15: 0] outgoing_data_to_and_from_the_cfi_flash_0;
  wire    [ 21: 0] p1_address_to_the_cfi_flash_0;
  wire    [  1: 0] p1_cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register;
  wire    [  1: 0] p1_cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register;
  wire             p1_read_n_to_the_cfi_flash_0;
  wire             p1_select_n_to_the_cfi_flash_0;
  wire             p1_write_n_to_the_cfi_flash_0;
  reg              read_n_to_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  reg              select_n_to_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  wire             time_to_write;
  wire             tri_state_bridge_0_avalon_slave_allgrants;
  wire             tri_state_bridge_0_avalon_slave_allow_new_arb_cycle;
  wire             tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant;
  wire             tri_state_bridge_0_avalon_slave_any_continuerequest;
  reg     [  1: 0] tri_state_bridge_0_avalon_slave_arb_addend;
  wire             tri_state_bridge_0_avalon_slave_arb_counter_enable;
  reg     [  1: 0] tri_state_bridge_0_avalon_slave_arb_share_counter;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_arb_share_counter_next_value;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_arb_share_set_values;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_arb_winner;
  wire             tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal;
  wire             tri_state_bridge_0_avalon_slave_beginbursttransfer_internal;
  wire             tri_state_bridge_0_avalon_slave_begins_xfer;
  wire    [  3: 0] tri_state_bridge_0_avalon_slave_chosen_master_double_vector;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_chosen_master_rot_left;
  wire             tri_state_bridge_0_avalon_slave_end_xfer;
  wire             tri_state_bridge_0_avalon_slave_firsttransfer;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_grant_vector;
  wire    [  1: 0] tri_state_bridge_0_avalon_slave_master_qreq_vector;
  wire             tri_state_bridge_0_avalon_slave_non_bursting_master_requests;
  wire             tri_state_bridge_0_avalon_slave_read_pending;
  reg              tri_state_bridge_0_avalon_slave_reg_firsttransfer;
  reg     [  1: 0] tri_state_bridge_0_avalon_slave_saved_chosen_master_vector;
  reg              tri_state_bridge_0_avalon_slave_slavearbiterlockenable;
  wire             tri_state_bridge_0_avalon_slave_slavearbiterlockenable2;
  wire             tri_state_bridge_0_avalon_slave_unreg_firsttransfer;
  wire             tri_state_bridge_0_avalon_slave_write_pending;
  wire             wait_for_cfi_flash_0_s1_counter;
  reg              write_n_to_the_cfi_flash_0 /* synthesis ALTERA_ATTRIBUTE = "FAST_OUTPUT_REGISTER=ON"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_reasons_to_wait <= 0;
      else 
        d1_reasons_to_wait <= ~tri_state_bridge_0_avalon_slave_end_xfer;
    end


  assign tri_state_bridge_0_avalon_slave_begins_xfer = ~d1_reasons_to_wait & ((cpu_0_data_master_qualified_request_cfi_flash_0_s1 | cpu_0_instruction_master_qualified_request_cfi_flash_0_s1));
  assign cpu_0_data_master_requests_cfi_flash_0_s1 = ({cpu_0_data_master_address_to_slave[24 : 22] , 22'b0} == 25'h1400000) & (cpu_0_data_master_read | cpu_0_data_master_write);
  //~select_n_to_the_cfi_flash_0 of type chipselect to ~p1_select_n_to_the_cfi_flash_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          select_n_to_the_cfi_flash_0 <= ~0;
      else 
        select_n_to_the_cfi_flash_0 <= p1_select_n_to_the_cfi_flash_0;
    end


  assign tri_state_bridge_0_avalon_slave_write_pending = 0;
  //tri_state_bridge_0/avalon_slave read pending calc, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_read_pending = 0;

  //tri_state_bridge_0_avalon_slave_arb_share_counter set values, which is an e_mux
  assign tri_state_bridge_0_avalon_slave_arb_share_set_values = (cpu_0_data_master_granted_cfi_flash_0_s1)? 2 :
    (cpu_0_instruction_master_granted_cfi_flash_0_s1)? 2 :
    (cpu_0_data_master_granted_cfi_flash_0_s1)? 2 :
    (cpu_0_instruction_master_granted_cfi_flash_0_s1)? 2 :
    1;

  //tri_state_bridge_0_avalon_slave_non_bursting_master_requests mux, which is an e_mux
  assign tri_state_bridge_0_avalon_slave_non_bursting_master_requests = cpu_0_data_master_requests_cfi_flash_0_s1 |
    cpu_0_instruction_master_requests_cfi_flash_0_s1 |
    cpu_0_data_master_requests_cfi_flash_0_s1 |
    cpu_0_instruction_master_requests_cfi_flash_0_s1;

  //tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant mux, which is an e_mux
  assign tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant = 0;

  //tri_state_bridge_0_avalon_slave_arb_share_counter_next_value assignment, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_arb_share_counter_next_value = tri_state_bridge_0_avalon_slave_firsttransfer ? (tri_state_bridge_0_avalon_slave_arb_share_set_values - 1) : |tri_state_bridge_0_avalon_slave_arb_share_counter ? (tri_state_bridge_0_avalon_slave_arb_share_counter - 1) : 0;

  //tri_state_bridge_0_avalon_slave_allgrants all slave grants, which is an e_mux
  assign tri_state_bridge_0_avalon_slave_allgrants = (|tri_state_bridge_0_avalon_slave_grant_vector) |
    (|tri_state_bridge_0_avalon_slave_grant_vector) |
    (|tri_state_bridge_0_avalon_slave_grant_vector) |
    (|tri_state_bridge_0_avalon_slave_grant_vector);

  //tri_state_bridge_0_avalon_slave_end_xfer assignment, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_end_xfer = ~(cfi_flash_0_s1_waits_for_read | cfi_flash_0_s1_waits_for_write);

  //end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave arb share counter enable term, which is an e_assign
  assign end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave = tri_state_bridge_0_avalon_slave_end_xfer & (~tri_state_bridge_0_avalon_slave_any_bursting_master_saved_grant | in_a_read_cycle | in_a_write_cycle);

  //tri_state_bridge_0_avalon_slave_arb_share_counter arbitration counter enable, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_arb_counter_enable = (end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave & tri_state_bridge_0_avalon_slave_allgrants) | (end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave & ~tri_state_bridge_0_avalon_slave_non_bursting_master_requests);

  //tri_state_bridge_0_avalon_slave_arb_share_counter counter, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tri_state_bridge_0_avalon_slave_arb_share_counter <= 0;
      else if (tri_state_bridge_0_avalon_slave_arb_counter_enable)
          tri_state_bridge_0_avalon_slave_arb_share_counter <= tri_state_bridge_0_avalon_slave_arb_share_counter_next_value;
    end


  //tri_state_bridge_0_avalon_slave_slavearbiterlockenable slave enables arbiterlock, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tri_state_bridge_0_avalon_slave_slavearbiterlockenable <= 0;
      else if ((|tri_state_bridge_0_avalon_slave_master_qreq_vector & end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave) | (end_xfer_arb_share_counter_term_tri_state_bridge_0_avalon_slave & ~tri_state_bridge_0_avalon_slave_non_bursting_master_requests))
          tri_state_bridge_0_avalon_slave_slavearbiterlockenable <= |tri_state_bridge_0_avalon_slave_arb_share_counter_next_value;
    end


  //cpu_0/data_master tri_state_bridge_0/avalon_slave arbiterlock, which is an e_assign
  assign cpu_0_data_master_arbiterlock = tri_state_bridge_0_avalon_slave_slavearbiterlockenable & cpu_0_data_master_continuerequest;

  //tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 slave enables arbiterlock2, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 = |tri_state_bridge_0_avalon_slave_arb_share_counter_next_value;

  //cpu_0/data_master tri_state_bridge_0/avalon_slave arbiterlock2, which is an e_assign
  assign cpu_0_data_master_arbiterlock2 = tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 & cpu_0_data_master_continuerequest;

  //cpu_0/instruction_master tri_state_bridge_0/avalon_slave arbiterlock, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock = tri_state_bridge_0_avalon_slave_slavearbiterlockenable & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master tri_state_bridge_0/avalon_slave arbiterlock2, which is an e_assign
  assign cpu_0_instruction_master_arbiterlock2 = tri_state_bridge_0_avalon_slave_slavearbiterlockenable2 & cpu_0_instruction_master_continuerequest;

  //cpu_0/instruction_master granted cfi_flash_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_instruction_master_granted_slave_cfi_flash_0_s1 <= 0;
      else 
        last_cycle_cpu_0_instruction_master_granted_slave_cfi_flash_0_s1 <= cpu_0_instruction_master_saved_grant_cfi_flash_0_s1 ? 1 : (tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal | ~cpu_0_instruction_master_requests_cfi_flash_0_s1) ? 0 : last_cycle_cpu_0_instruction_master_granted_slave_cfi_flash_0_s1;
    end


  //cpu_0_instruction_master_continuerequest continued request, which is an e_mux
  assign cpu_0_instruction_master_continuerequest = last_cycle_cpu_0_instruction_master_granted_slave_cfi_flash_0_s1 & cpu_0_instruction_master_requests_cfi_flash_0_s1;

  //tri_state_bridge_0_avalon_slave_any_continuerequest at least one master continues requesting, which is an e_mux
  assign tri_state_bridge_0_avalon_slave_any_continuerequest = cpu_0_instruction_master_continuerequest |
    cpu_0_data_master_continuerequest;

  assign cpu_0_data_master_qualified_request_cfi_flash_0_s1 = cpu_0_data_master_requests_cfi_flash_0_s1 & ~((cpu_0_data_master_read & (tri_state_bridge_0_avalon_slave_write_pending | (tri_state_bridge_0_avalon_slave_read_pending) | (2 < cpu_0_data_master_latency_counter) | (|cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register))) | ((tri_state_bridge_0_avalon_slave_read_pending | !cpu_0_data_master_byteenable_cfi_flash_0_s1) & cpu_0_data_master_write) | cpu_0_instruction_master_arbiterlock);
  //cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in = cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_read & ~cfi_flash_0_s1_waits_for_read;

  //shift register p1 cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register = {cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register, cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register_in};

  //cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register <= 0;
      else 
        cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register <= p1_cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register;
    end


  //local readdatavalid cpu_0_data_master_read_data_valid_cfi_flash_0_s1, which is an e_mux
  assign cpu_0_data_master_read_data_valid_cfi_flash_0_s1 = cpu_0_data_master_read_data_valid_cfi_flash_0_s1_shift_register[1];

  //data_to_and_from_the_cfi_flash_0 register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          incoming_data_to_and_from_the_cfi_flash_0 <= 0;
      else 
        incoming_data_to_and_from_the_cfi_flash_0 <= data_to_and_from_the_cfi_flash_0;
    end


  //cfi_flash_0_s1_with_write_latency assignment, which is an e_assign
  assign cfi_flash_0_s1_with_write_latency = in_a_write_cycle & (cpu_0_data_master_qualified_request_cfi_flash_0_s1 | cpu_0_instruction_master_qualified_request_cfi_flash_0_s1);

  //time to write the data, which is an e_mux
  assign time_to_write = (cfi_flash_0_s1_with_write_latency)? 1 :
    0;

  //d1_outgoing_data_to_and_from_the_cfi_flash_0 register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_outgoing_data_to_and_from_the_cfi_flash_0 <= 0;
      else 
        d1_outgoing_data_to_and_from_the_cfi_flash_0 <= outgoing_data_to_and_from_the_cfi_flash_0;
    end


  //write cycle delayed by 1, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_in_a_write_cycle <= 0;
      else 
        d1_in_a_write_cycle <= time_to_write;
    end


  //d1_outgoing_data_to_and_from_the_cfi_flash_0 tristate driver, which is an e_assign
  assign data_to_and_from_the_cfi_flash_0 = (d1_in_a_write_cycle)? d1_outgoing_data_to_and_from_the_cfi_flash_0:{16{1'bz}};

  //outgoing_data_to_and_from_the_cfi_flash_0 mux, which is an e_mux
  assign outgoing_data_to_and_from_the_cfi_flash_0 = cpu_0_data_master_dbs_write_16;

  assign cpu_0_instruction_master_requests_cfi_flash_0_s1 = (({cpu_0_instruction_master_address_to_slave[24 : 22] , 22'b0} == 25'h1400000) & (cpu_0_instruction_master_read)) & cpu_0_instruction_master_read;
  //cpu_0/data_master granted cfi_flash_0/s1 last time, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          last_cycle_cpu_0_data_master_granted_slave_cfi_flash_0_s1 <= 0;
      else 
        last_cycle_cpu_0_data_master_granted_slave_cfi_flash_0_s1 <= cpu_0_data_master_saved_grant_cfi_flash_0_s1 ? 1 : (tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal | ~cpu_0_data_master_requests_cfi_flash_0_s1) ? 0 : last_cycle_cpu_0_data_master_granted_slave_cfi_flash_0_s1;
    end


  //cpu_0_data_master_continuerequest continued request, which is an e_mux
  assign cpu_0_data_master_continuerequest = last_cycle_cpu_0_data_master_granted_slave_cfi_flash_0_s1 & cpu_0_data_master_requests_cfi_flash_0_s1;

  assign cpu_0_instruction_master_qualified_request_cfi_flash_0_s1 = cpu_0_instruction_master_requests_cfi_flash_0_s1 & ~((cpu_0_instruction_master_read & (tri_state_bridge_0_avalon_slave_write_pending | (tri_state_bridge_0_avalon_slave_read_pending) | (2 < cpu_0_instruction_master_latency_counter) | (|cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register))) | cpu_0_data_master_arbiterlock);
  //cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in mux for readlatency shift register, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in = cpu_0_instruction_master_granted_cfi_flash_0_s1 & cpu_0_instruction_master_read & ~cfi_flash_0_s1_waits_for_read;

  //shift register p1 cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register in if flush, otherwise shift left, which is an e_mux
  assign p1_cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register = {cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register, cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register_in};

  //cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register for remembering which master asked for a fixed latency read, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register <= 0;
      else 
        cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register <= p1_cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register;
    end


  //local readdatavalid cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1, which is an e_mux
  assign cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1 = cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1_shift_register[1];

  //allow new arb cycle for tri_state_bridge_0/avalon_slave, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_allow_new_arb_cycle = ~cpu_0_data_master_arbiterlock & ~cpu_0_instruction_master_arbiterlock;

  //cpu_0/instruction_master assignment into master qualified-requests vector for cfi_flash_0/s1, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_master_qreq_vector[0] = cpu_0_instruction_master_qualified_request_cfi_flash_0_s1;

  //cpu_0/instruction_master grant cfi_flash_0/s1, which is an e_assign
  assign cpu_0_instruction_master_granted_cfi_flash_0_s1 = tri_state_bridge_0_avalon_slave_grant_vector[0];

  //cpu_0/instruction_master saved-grant cfi_flash_0/s1, which is an e_assign
  assign cpu_0_instruction_master_saved_grant_cfi_flash_0_s1 = tri_state_bridge_0_avalon_slave_arb_winner[0] && cpu_0_instruction_master_requests_cfi_flash_0_s1;

  //cpu_0/data_master assignment into master qualified-requests vector for cfi_flash_0/s1, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_master_qreq_vector[1] = cpu_0_data_master_qualified_request_cfi_flash_0_s1;

  //cpu_0/data_master grant cfi_flash_0/s1, which is an e_assign
  assign cpu_0_data_master_granted_cfi_flash_0_s1 = tri_state_bridge_0_avalon_slave_grant_vector[1];

  //cpu_0/data_master saved-grant cfi_flash_0/s1, which is an e_assign
  assign cpu_0_data_master_saved_grant_cfi_flash_0_s1 = tri_state_bridge_0_avalon_slave_arb_winner[1] && cpu_0_data_master_requests_cfi_flash_0_s1;

  //tri_state_bridge_0/avalon_slave chosen-master double-vector, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_chosen_master_double_vector = {tri_state_bridge_0_avalon_slave_master_qreq_vector, tri_state_bridge_0_avalon_slave_master_qreq_vector} & ({~tri_state_bridge_0_avalon_slave_master_qreq_vector, ~tri_state_bridge_0_avalon_slave_master_qreq_vector} + tri_state_bridge_0_avalon_slave_arb_addend);

  //stable onehot encoding of arb winner
  assign tri_state_bridge_0_avalon_slave_arb_winner = (tri_state_bridge_0_avalon_slave_allow_new_arb_cycle & | tri_state_bridge_0_avalon_slave_grant_vector) ? tri_state_bridge_0_avalon_slave_grant_vector : tri_state_bridge_0_avalon_slave_saved_chosen_master_vector;

  //saved tri_state_bridge_0_avalon_slave_grant_vector, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tri_state_bridge_0_avalon_slave_saved_chosen_master_vector <= 0;
      else if (tri_state_bridge_0_avalon_slave_allow_new_arb_cycle)
          tri_state_bridge_0_avalon_slave_saved_chosen_master_vector <= |tri_state_bridge_0_avalon_slave_grant_vector ? tri_state_bridge_0_avalon_slave_grant_vector : tri_state_bridge_0_avalon_slave_saved_chosen_master_vector;
    end


  //onehot encoding of chosen master
  assign tri_state_bridge_0_avalon_slave_grant_vector = {(tri_state_bridge_0_avalon_slave_chosen_master_double_vector[1] | tri_state_bridge_0_avalon_slave_chosen_master_double_vector[3]),
    (tri_state_bridge_0_avalon_slave_chosen_master_double_vector[0] | tri_state_bridge_0_avalon_slave_chosen_master_double_vector[2])};

  //tri_state_bridge_0/avalon_slave chosen master rotated left, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_chosen_master_rot_left = (tri_state_bridge_0_avalon_slave_arb_winner << 1) ? (tri_state_bridge_0_avalon_slave_arb_winner << 1) : 1;

  //tri_state_bridge_0/avalon_slave's addend for next-master-grant
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tri_state_bridge_0_avalon_slave_arb_addend <= 1;
      else if (|tri_state_bridge_0_avalon_slave_grant_vector)
          tri_state_bridge_0_avalon_slave_arb_addend <= tri_state_bridge_0_avalon_slave_end_xfer? tri_state_bridge_0_avalon_slave_chosen_master_rot_left : tri_state_bridge_0_avalon_slave_grant_vector;
    end


  assign p1_select_n_to_the_cfi_flash_0 = ~(cpu_0_data_master_granted_cfi_flash_0_s1 | cpu_0_instruction_master_granted_cfi_flash_0_s1);
  //tri_state_bridge_0_avalon_slave_firsttransfer first transaction, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_firsttransfer = tri_state_bridge_0_avalon_slave_begins_xfer ? tri_state_bridge_0_avalon_slave_unreg_firsttransfer : tri_state_bridge_0_avalon_slave_reg_firsttransfer;

  //tri_state_bridge_0_avalon_slave_unreg_firsttransfer first transaction, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_unreg_firsttransfer = ~(tri_state_bridge_0_avalon_slave_slavearbiterlockenable & tri_state_bridge_0_avalon_slave_any_continuerequest);

  //tri_state_bridge_0_avalon_slave_reg_firsttransfer first transaction, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          tri_state_bridge_0_avalon_slave_reg_firsttransfer <= 1'b1;
      else if (tri_state_bridge_0_avalon_slave_begins_xfer)
          tri_state_bridge_0_avalon_slave_reg_firsttransfer <= tri_state_bridge_0_avalon_slave_unreg_firsttransfer;
    end


  //tri_state_bridge_0_avalon_slave_beginbursttransfer_internal begin burst transfer, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_beginbursttransfer_internal = tri_state_bridge_0_avalon_slave_begins_xfer;

  //tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal arbitration_holdoff, which is an e_assign
  assign tri_state_bridge_0_avalon_slave_arbitration_holdoff_internal = tri_state_bridge_0_avalon_slave_begins_xfer & tri_state_bridge_0_avalon_slave_firsttransfer;

  //~read_n_to_the_cfi_flash_0 of type read to ~p1_read_n_to_the_cfi_flash_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          read_n_to_the_cfi_flash_0 <= ~0;
      else 
        read_n_to_the_cfi_flash_0 <= p1_read_n_to_the_cfi_flash_0;
    end


  //~p1_read_n_to_the_cfi_flash_0 assignment, which is an e_mux
  assign p1_read_n_to_the_cfi_flash_0 = ~(((cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_cfi_flash_0_s1 & cpu_0_instruction_master_read))& ~tri_state_bridge_0_avalon_slave_begins_xfer & (cfi_flash_0_s1_wait_counter < 8));

  //~write_n_to_the_cfi_flash_0 of type write to ~p1_write_n_to_the_cfi_flash_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          write_n_to_the_cfi_flash_0 <= ~0;
      else 
        write_n_to_the_cfi_flash_0 <= p1_write_n_to_the_cfi_flash_0;
    end


  //~p1_write_n_to_the_cfi_flash_0 assignment, which is an e_mux
  assign p1_write_n_to_the_cfi_flash_0 = ~(((cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_write)) & ~tri_state_bridge_0_avalon_slave_begins_xfer & (cfi_flash_0_s1_wait_counter >= 2) & (cfi_flash_0_s1_wait_counter < 10));

  //address_to_the_cfi_flash_0 of type address to p1_address_to_the_cfi_flash_0, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          address_to_the_cfi_flash_0 <= 0;
      else 
        address_to_the_cfi_flash_0 <= p1_address_to_the_cfi_flash_0;
    end


  //p1_address_to_the_cfi_flash_0 mux, which is an e_mux
  assign p1_address_to_the_cfi_flash_0 = (cpu_0_data_master_granted_cfi_flash_0_s1)? ({cpu_0_data_master_address_to_slave >> 2,
    cpu_0_data_master_dbs_address[1],
    {1 {1'b0}}}) :
    ({cpu_0_instruction_master_address_to_slave >> 2,
    cpu_0_instruction_master_dbs_address[1],
    {1 {1'b0}}});

  //d1_tri_state_bridge_0_avalon_slave_end_xfer register, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          d1_tri_state_bridge_0_avalon_slave_end_xfer <= 1;
      else 
        d1_tri_state_bridge_0_avalon_slave_end_xfer <= tri_state_bridge_0_avalon_slave_end_xfer;
    end


  //cfi_flash_0_s1_waits_for_read in a cycle, which is an e_mux
  assign cfi_flash_0_s1_waits_for_read = cfi_flash_0_s1_in_a_read_cycle & wait_for_cfi_flash_0_s1_counter;

  //cfi_flash_0_s1_in_a_read_cycle assignment, which is an e_assign
  assign cfi_flash_0_s1_in_a_read_cycle = (cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_read) | (cpu_0_instruction_master_granted_cfi_flash_0_s1 & cpu_0_instruction_master_read);

  //in_a_read_cycle assignment, which is an e_mux
  assign in_a_read_cycle = cfi_flash_0_s1_in_a_read_cycle;

  //cfi_flash_0_s1_waits_for_write in a cycle, which is an e_mux
  assign cfi_flash_0_s1_waits_for_write = cfi_flash_0_s1_in_a_write_cycle & wait_for_cfi_flash_0_s1_counter;

  //cfi_flash_0_s1_in_a_write_cycle assignment, which is an e_assign
  assign cfi_flash_0_s1_in_a_write_cycle = cpu_0_data_master_granted_cfi_flash_0_s1 & cpu_0_data_master_write;

  //in_a_write_cycle assignment, which is an e_mux
  assign in_a_write_cycle = cfi_flash_0_s1_in_a_write_cycle;

  assign cfi_flash_0_s1_wait_counter_eq_0 = cfi_flash_0_s1_wait_counter == 0;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          cfi_flash_0_s1_wait_counter <= 0;
      else 
        cfi_flash_0_s1_wait_counter <= cfi_flash_0_s1_counter_load_value;
    end


  assign cfi_flash_0_s1_counter_load_value = ((cfi_flash_0_s1_in_a_write_cycle & tri_state_bridge_0_avalon_slave_begins_xfer))? 10 :
    ((cfi_flash_0_s1_in_a_read_cycle & tri_state_bridge_0_avalon_slave_begins_xfer))? 8 :
    (~cfi_flash_0_s1_wait_counter_eq_0)? cfi_flash_0_s1_wait_counter - 1 :
    0;

  assign wait_for_cfi_flash_0_s1_counter = tri_state_bridge_0_avalon_slave_begins_xfer | ~cfi_flash_0_s1_wait_counter_eq_0;
  assign {cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_1,
cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_0} = cpu_0_data_master_byteenable;
  assign cpu_0_data_master_byteenable_cfi_flash_0_s1 = ((cpu_0_data_master_dbs_address[1] == 0))? cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_0 :
    cpu_0_data_master_byteenable_cfi_flash_0_s1_segment_1;


//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  //incoming_data_to_and_from_the_cfi_flash_0_bit_0_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_0_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[0]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[0] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[0] = incoming_data_to_and_from_the_cfi_flash_0_bit_0_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[0];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_1_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_1_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[1]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[1] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[1] = incoming_data_to_and_from_the_cfi_flash_0_bit_1_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[1];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_2_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_2_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[2]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[2] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[2] = incoming_data_to_and_from_the_cfi_flash_0_bit_2_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[2];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_3_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_3_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[3]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[3] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[3] = incoming_data_to_and_from_the_cfi_flash_0_bit_3_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[3];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_4_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_4_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[4]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[4] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[4] = incoming_data_to_and_from_the_cfi_flash_0_bit_4_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[4];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_5_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_5_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[5]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[5] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[5] = incoming_data_to_and_from_the_cfi_flash_0_bit_5_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[5];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_6_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_6_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[6]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[6] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[6] = incoming_data_to_and_from_the_cfi_flash_0_bit_6_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[6];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_7_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_7_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[7]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[7] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[7] = incoming_data_to_and_from_the_cfi_flash_0_bit_7_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[7];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_8_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_8_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[8]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[8] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[8] = incoming_data_to_and_from_the_cfi_flash_0_bit_8_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[8];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_9_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_9_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[9]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[9] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[9] = incoming_data_to_and_from_the_cfi_flash_0_bit_9_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[9];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_10_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_10_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[10]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[10] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[10] = incoming_data_to_and_from_the_cfi_flash_0_bit_10_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[10];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_11_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_11_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[11]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[11] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[11] = incoming_data_to_and_from_the_cfi_flash_0_bit_11_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[11];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_12_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_12_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[12]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[12] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[12] = incoming_data_to_and_from_the_cfi_flash_0_bit_12_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[12];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_13_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_13_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[13]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[13] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[13] = incoming_data_to_and_from_the_cfi_flash_0_bit_13_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[13];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_14_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_14_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[14]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[14] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[14] = incoming_data_to_and_from_the_cfi_flash_0_bit_14_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[14];

  //incoming_data_to_and_from_the_cfi_flash_0_bit_15_is_x x check, which is an e_assign_is_x
  assign incoming_data_to_and_from_the_cfi_flash_0_bit_15_is_x = ^(incoming_data_to_and_from_the_cfi_flash_0[15]) === 1'bx;

  //Crush incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[15] Xs to 0, which is an e_assign
  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0[15] = incoming_data_to_and_from_the_cfi_flash_0_bit_15_is_x ? 1'b0 : incoming_data_to_and_from_the_cfi_flash_0[15];

  //cfi_flash_0/s1 enable non-zero assertions, which is an e_register
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          enable_nonzero_assertions <= 0;
      else 
        enable_nonzero_assertions <= 1'b1;
    end


  //grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_granted_cfi_flash_0_s1 + cpu_0_instruction_master_granted_cfi_flash_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of grant signals are active simultaneously", $time);
          $stop;
        end
    end


  //saved_grant signals are active simultaneously, which is an e_process
  always @(posedge clk)
    begin
      if (cpu_0_data_master_saved_grant_cfi_flash_0_s1 + cpu_0_instruction_master_saved_grant_cfi_flash_0_s1 > 1)
        begin
          $write("%0d ns: > 1 of saved_grant signals are active simultaneously", $time);
          $stop;
        end
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  
//  assign incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0 = incoming_data_to_and_from_the_cfi_flash_0;
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module tri_state_bridge_0_bridge_arbitrator 
;



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nioscpu_reset_clk_0_domain_synch_module (
                                                 // inputs:
                                                  clk,
                                                  data_in,
                                                  reset_n,

                                                 // outputs:
                                                  data_out
                                               )
;

  output           data_out;
  input            clk;
  input            data_in;
  input            reset_n;

  reg              data_in_d1 /* synthesis ALTERA_ATTRIBUTE = "{-from \"*\"} CUT=ON ; PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  reg              data_out /* synthesis ALTERA_ATTRIBUTE = "PRESERVE_REGISTER=ON ; SUPPRESS_DA_RULE_INTERNAL=R101"  */;
  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_in_d1 <= 0;
      else 
        data_in_d1 <= data_in;
    end


  always @(posedge clk or negedge reset_n)
    begin
      if (reset_n == 0)
          data_out <= 0;
      else 
        data_out <= data_in_d1;
    end



endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module nioscpu (
                 // 1) global signals:
                  clk_0,
                  reset_n,

                 // the_button_pio
                  in_port_to_the_button_pio,

                 // the_col
                  out_port_from_the_col,

                 // the_led_pio
                  out_port_from_the_led_pio,

                 // the_row
                  out_port_from_the_row,

                 // the_sdram_0
                  zs_addr_from_the_sdram_0,
                  zs_ba_from_the_sdram_0,
                  zs_cas_n_from_the_sdram_0,
                  zs_cke_from_the_sdram_0,
                  zs_cs_n_from_the_sdram_0,
                  zs_dq_to_and_from_the_sdram_0,
                  zs_dqm_from_the_sdram_0,
                  zs_ras_n_from_the_sdram_0,
                  zs_we_n_from_the_sdram_0,

                 // the_tft_lcd_data
                  out_port_from_the_tft_lcd_data,

                 // the_tft_lcd_nrd
                  out_port_from_the_tft_lcd_nrd,

                 // the_tft_lcd_nrst
                  out_port_from_the_tft_lcd_nrst,

                 // the_tft_lcd_nwr
                  out_port_from_the_tft_lcd_nwr,

                 // the_tft_lcd_rs
                  out_port_from_the_tft_lcd_rs,

                 // the_tri_state_bridge_0_avalon_slave
                  address_to_the_cfi_flash_0,
                  data_to_and_from_the_cfi_flash_0,
                  read_n_to_the_cfi_flash_0,
                  select_n_to_the_cfi_flash_0,
                  write_n_to_the_cfi_flash_0
               )
;

  output  [ 21: 0] address_to_the_cfi_flash_0;
  inout   [ 15: 0] data_to_and_from_the_cfi_flash_0;
  output  [  3: 0] out_port_from_the_col;
  output  [  7: 0] out_port_from_the_led_pio;
  output  [ 15: 0] out_port_from_the_row;
  output  [  7: 0] out_port_from_the_tft_lcd_data;
  output           out_port_from_the_tft_lcd_nrd;
  output           out_port_from_the_tft_lcd_nrst;
  output           out_port_from_the_tft_lcd_nwr;
  output           out_port_from_the_tft_lcd_rs;
  output           read_n_to_the_cfi_flash_0;
  output           select_n_to_the_cfi_flash_0;
  output           write_n_to_the_cfi_flash_0;
  output  [ 11: 0] zs_addr_from_the_sdram_0;
  output  [  1: 0] zs_ba_from_the_sdram_0;
  output           zs_cas_n_from_the_sdram_0;
  output           zs_cke_from_the_sdram_0;
  output           zs_cs_n_from_the_sdram_0;
  inout   [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  output  [  1: 0] zs_dqm_from_the_sdram_0;
  output           zs_ras_n_from_the_sdram_0;
  output           zs_we_n_from_the_sdram_0;
  input            clk_0;
  input   [  7: 0] in_port_to_the_button_pio;
  input            reset_n;

  wire    [ 21: 0] address_to_the_cfi_flash_0;
  wire    [  1: 0] button_pio_s1_address;
  wire             button_pio_s1_chipselect;
  wire             button_pio_s1_irq;
  wire             button_pio_s1_irq_from_sa;
  wire    [  7: 0] button_pio_s1_readdata;
  wire    [  7: 0] button_pio_s1_readdata_from_sa;
  wire             button_pio_s1_reset_n;
  wire             button_pio_s1_write_n;
  wire    [  7: 0] button_pio_s1_writedata;
  wire             cfi_flash_0_s1_wait_counter_eq_0;
  wire             clk_0_reset_n;
  wire    [  1: 0] col_s1_address;
  wire             col_s1_chipselect;
  wire    [  3: 0] col_s1_readdata;
  wire    [  3: 0] col_s1_readdata_from_sa;
  wire             col_s1_reset_n;
  wire             col_s1_write_n;
  wire    [  3: 0] col_s1_writedata;
  wire    [ 24: 0] cpu_0_data_master_address;
  wire    [ 24: 0] cpu_0_data_master_address_to_slave;
  wire    [  3: 0] cpu_0_data_master_byteenable;
  wire    [  1: 0] cpu_0_data_master_byteenable_cfi_flash_0_s1;
  wire    [  1: 0] cpu_0_data_master_byteenable_sdram_0_s1;
  wire    [  1: 0] cpu_0_data_master_dbs_address;
  wire    [ 15: 0] cpu_0_data_master_dbs_write_16;
  wire             cpu_0_data_master_debugaccess;
  wire             cpu_0_data_master_granted_button_pio_s1;
  wire             cpu_0_data_master_granted_cfi_flash_0_s1;
  wire             cpu_0_data_master_granted_col_s1;
  wire             cpu_0_data_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_granted_led_pio_s1;
  wire             cpu_0_data_master_granted_row_s1;
  wire             cpu_0_data_master_granted_sdram_0_s1;
  wire             cpu_0_data_master_granted_tft_lcd_data_s1;
  wire             cpu_0_data_master_granted_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_granted_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_granted_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_granted_tft_lcd_rs_s1;
  wire    [ 31: 0] cpu_0_data_master_irq;
  wire    [  1: 0] cpu_0_data_master_latency_counter;
  wire             cpu_0_data_master_qualified_request_button_pio_s1;
  wire             cpu_0_data_master_qualified_request_cfi_flash_0_s1;
  wire             cpu_0_data_master_qualified_request_col_s1;
  wire             cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_qualified_request_led_pio_s1;
  wire             cpu_0_data_master_qualified_request_row_s1;
  wire             cpu_0_data_master_qualified_request_sdram_0_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_data_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_qualified_request_tft_lcd_rs_s1;
  wire             cpu_0_data_master_read;
  wire             cpu_0_data_master_read_data_valid_button_pio_s1;
  wire             cpu_0_data_master_read_data_valid_cfi_flash_0_s1;
  wire             cpu_0_data_master_read_data_valid_col_s1;
  wire             cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_read_data_valid_led_pio_s1;
  wire             cpu_0_data_master_read_data_valid_row_s1;
  wire             cpu_0_data_master_read_data_valid_sdram_0_s1;
  wire             cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_data_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_read_data_valid_tft_lcd_rs_s1;
  wire    [ 31: 0] cpu_0_data_master_readdata;
  wire             cpu_0_data_master_readdatavalid;
  wire             cpu_0_data_master_requests_button_pio_s1;
  wire             cpu_0_data_master_requests_cfi_flash_0_s1;
  wire             cpu_0_data_master_requests_col_s1;
  wire             cpu_0_data_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave;
  wire             cpu_0_data_master_requests_led_pio_s1;
  wire             cpu_0_data_master_requests_row_s1;
  wire             cpu_0_data_master_requests_sdram_0_s1;
  wire             cpu_0_data_master_requests_tft_lcd_data_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nrd_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nrst_s1;
  wire             cpu_0_data_master_requests_tft_lcd_nwr_s1;
  wire             cpu_0_data_master_requests_tft_lcd_rs_s1;
  wire             cpu_0_data_master_waitrequest;
  wire             cpu_0_data_master_write;
  wire    [ 31: 0] cpu_0_data_master_writedata;
  wire    [ 24: 0] cpu_0_instruction_master_address;
  wire    [ 24: 0] cpu_0_instruction_master_address_to_slave;
  wire    [  1: 0] cpu_0_instruction_master_dbs_address;
  wire             cpu_0_instruction_master_granted_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_granted_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_granted_sdram_0_s1;
  wire             cpu_0_instruction_master_granted_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_granted_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_granted_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_granted_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_granted_tft_lcd_rs_s1;
  wire    [  1: 0] cpu_0_instruction_master_latency_counter;
  wire             cpu_0_instruction_master_qualified_request_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_qualified_request_sdram_0_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_read;
  wire             cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_read_data_valid_sdram_0_s1;
  wire             cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1;
  wire    [ 31: 0] cpu_0_instruction_master_readdata;
  wire             cpu_0_instruction_master_readdatavalid;
  wire             cpu_0_instruction_master_requests_cfi_flash_0_s1;
  wire             cpu_0_instruction_master_requests_cpu_0_jtag_debug_module;
  wire             cpu_0_instruction_master_requests_sdram_0_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_data_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nrd_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nrst_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_nwr_s1;
  wire             cpu_0_instruction_master_requests_tft_lcd_rs_s1;
  wire             cpu_0_instruction_master_waitrequest;
  wire    [  8: 0] cpu_0_jtag_debug_module_address;
  wire             cpu_0_jtag_debug_module_begintransfer;
  wire    [  3: 0] cpu_0_jtag_debug_module_byteenable;
  wire             cpu_0_jtag_debug_module_chipselect;
  wire             cpu_0_jtag_debug_module_debugaccess;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata;
  wire    [ 31: 0] cpu_0_jtag_debug_module_readdata_from_sa;
  wire             cpu_0_jtag_debug_module_reset;
  wire             cpu_0_jtag_debug_module_reset_n;
  wire             cpu_0_jtag_debug_module_resetrequest;
  wire             cpu_0_jtag_debug_module_resetrequest_from_sa;
  wire             cpu_0_jtag_debug_module_write;
  wire    [ 31: 0] cpu_0_jtag_debug_module_writedata;
  wire             d1_button_pio_s1_end_xfer;
  wire             d1_col_s1_end_xfer;
  wire             d1_cpu_0_jtag_debug_module_end_xfer;
  wire             d1_jtag_uart_0_avalon_jtag_slave_end_xfer;
  wire             d1_led_pio_s1_end_xfer;
  wire             d1_row_s1_end_xfer;
  wire             d1_sdram_0_s1_end_xfer;
  wire             d1_tft_lcd_data_s1_end_xfer;
  wire             d1_tft_lcd_nrd_s1_end_xfer;
  wire             d1_tft_lcd_nrst_s1_end_xfer;
  wire             d1_tft_lcd_nwr_s1_end_xfer;
  wire             d1_tft_lcd_rs_s1_end_xfer;
  wire             d1_tri_state_bridge_0_avalon_slave_end_xfer;
  wire    [ 15: 0] data_to_and_from_the_cfi_flash_0;
  wire    [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0;
  wire    [ 15: 0] incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0;
  wire             jtag_uart_0_avalon_jtag_slave_address;
  wire             jtag_uart_0_avalon_jtag_slave_chipselect;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_irq;
  wire             jtag_uart_0_avalon_jtag_slave_irq_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_read_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_readdata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_reset_n;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest;
  wire             jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_write_n;
  wire    [ 31: 0] jtag_uart_0_avalon_jtag_slave_writedata;
  wire    [  1: 0] led_pio_s1_address;
  wire             led_pio_s1_chipselect;
  wire    [  7: 0] led_pio_s1_readdata;
  wire    [  7: 0] led_pio_s1_readdata_from_sa;
  wire             led_pio_s1_reset_n;
  wire             led_pio_s1_write_n;
  wire    [  7: 0] led_pio_s1_writedata;
  wire    [  3: 0] out_port_from_the_col;
  wire    [  7: 0] out_port_from_the_led_pio;
  wire    [ 15: 0] out_port_from_the_row;
  wire    [  7: 0] out_port_from_the_tft_lcd_data;
  wire             out_port_from_the_tft_lcd_nrd;
  wire             out_port_from_the_tft_lcd_nrst;
  wire             out_port_from_the_tft_lcd_nwr;
  wire             out_port_from_the_tft_lcd_rs;
  wire             read_n_to_the_cfi_flash_0;
  wire             reset_n_sources;
  wire    [  1: 0] row_s1_address;
  wire             row_s1_chipselect;
  wire    [ 15: 0] row_s1_readdata;
  wire    [ 15: 0] row_s1_readdata_from_sa;
  wire             row_s1_reset_n;
  wire             row_s1_write_n;
  wire    [ 15: 0] row_s1_writedata;
  wire    [ 21: 0] sdram_0_s1_address;
  wire    [  1: 0] sdram_0_s1_byteenable_n;
  wire             sdram_0_s1_chipselect;
  wire             sdram_0_s1_read_n;
  wire    [ 15: 0] sdram_0_s1_readdata;
  wire    [ 15: 0] sdram_0_s1_readdata_from_sa;
  wire             sdram_0_s1_readdatavalid;
  wire             sdram_0_s1_reset_n;
  wire             sdram_0_s1_waitrequest;
  wire             sdram_0_s1_waitrequest_from_sa;
  wire             sdram_0_s1_write_n;
  wire    [ 15: 0] sdram_0_s1_writedata;
  wire             select_n_to_the_cfi_flash_0;
  wire    [  1: 0] tft_lcd_data_s1_address;
  wire             tft_lcd_data_s1_chipselect;
  wire    [  7: 0] tft_lcd_data_s1_readdata;
  wire    [  7: 0] tft_lcd_data_s1_readdata_from_sa;
  wire             tft_lcd_data_s1_reset_n;
  wire             tft_lcd_data_s1_write_n;
  wire    [  7: 0] tft_lcd_data_s1_writedata;
  wire    [  1: 0] tft_lcd_nrd_s1_address;
  wire             tft_lcd_nrd_s1_chipselect;
  wire             tft_lcd_nrd_s1_readdata;
  wire             tft_lcd_nrd_s1_readdata_from_sa;
  wire             tft_lcd_nrd_s1_reset_n;
  wire             tft_lcd_nrd_s1_write_n;
  wire             tft_lcd_nrd_s1_writedata;
  wire    [  1: 0] tft_lcd_nrst_s1_address;
  wire             tft_lcd_nrst_s1_chipselect;
  wire             tft_lcd_nrst_s1_readdata;
  wire             tft_lcd_nrst_s1_readdata_from_sa;
  wire             tft_lcd_nrst_s1_reset_n;
  wire             tft_lcd_nrst_s1_write_n;
  wire             tft_lcd_nrst_s1_writedata;
  wire    [  1: 0] tft_lcd_nwr_s1_address;
  wire             tft_lcd_nwr_s1_chipselect;
  wire             tft_lcd_nwr_s1_readdata;
  wire             tft_lcd_nwr_s1_readdata_from_sa;
  wire             tft_lcd_nwr_s1_reset_n;
  wire             tft_lcd_nwr_s1_write_n;
  wire             tft_lcd_nwr_s1_writedata;
  wire    [  1: 0] tft_lcd_rs_s1_address;
  wire             tft_lcd_rs_s1_chipselect;
  wire             tft_lcd_rs_s1_readdata;
  wire             tft_lcd_rs_s1_readdata_from_sa;
  wire             tft_lcd_rs_s1_reset_n;
  wire             tft_lcd_rs_s1_write_n;
  wire             tft_lcd_rs_s1_writedata;
  wire             write_n_to_the_cfi_flash_0;
  wire    [ 11: 0] zs_addr_from_the_sdram_0;
  wire    [  1: 0] zs_ba_from_the_sdram_0;
  wire             zs_cas_n_from_the_sdram_0;
  wire             zs_cke_from_the_sdram_0;
  wire             zs_cs_n_from_the_sdram_0;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  wire    [  1: 0] zs_dqm_from_the_sdram_0;
  wire             zs_ras_n_from_the_sdram_0;
  wire             zs_we_n_from_the_sdram_0;
  button_pio_s1_arbitrator the_button_pio_s1
    (
      .button_pio_s1_address                                       (button_pio_s1_address),
      .button_pio_s1_chipselect                                    (button_pio_s1_chipselect),
      .button_pio_s1_irq                                           (button_pio_s1_irq),
      .button_pio_s1_irq_from_sa                                   (button_pio_s1_irq_from_sa),
      .button_pio_s1_readdata                                      (button_pio_s1_readdata),
      .button_pio_s1_readdata_from_sa                              (button_pio_s1_readdata_from_sa),
      .button_pio_s1_reset_n                                       (button_pio_s1_reset_n),
      .button_pio_s1_write_n                                       (button_pio_s1_write_n),
      .button_pio_s1_writedata                                     (button_pio_s1_writedata),
      .clk                                                         (clk_0),
      .cpu_0_data_master_address_to_slave                          (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_button_pio_s1                     (cpu_0_data_master_granted_button_pio_s1),
      .cpu_0_data_master_latency_counter                           (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_button_pio_s1           (cpu_0_data_master_qualified_request_button_pio_s1),
      .cpu_0_data_master_read                                      (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_button_pio_s1             (cpu_0_data_master_read_data_valid_button_pio_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_button_pio_s1                    (cpu_0_data_master_requests_button_pio_s1),
      .cpu_0_data_master_write                                     (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                 (cpu_0_data_master_writedata),
      .d1_button_pio_s1_end_xfer                                   (d1_button_pio_s1_end_xfer),
      .reset_n                                                     (clk_0_reset_n)
    );

  button_pio the_button_pio
    (
      .address    (button_pio_s1_address),
      .chipselect (button_pio_s1_chipselect),
      .clk        (clk_0),
      .in_port    (in_port_to_the_button_pio),
      .irq        (button_pio_s1_irq),
      .readdata   (button_pio_s1_readdata),
      .reset_n    (button_pio_s1_reset_n),
      .write_n    (button_pio_s1_write_n),
      .writedata  (button_pio_s1_writedata)
    );

  col_s1_arbitrator the_col_s1
    (
      .clk                                                         (clk_0),
      .col_s1_address                                              (col_s1_address),
      .col_s1_chipselect                                           (col_s1_chipselect),
      .col_s1_readdata                                             (col_s1_readdata),
      .col_s1_readdata_from_sa                                     (col_s1_readdata_from_sa),
      .col_s1_reset_n                                              (col_s1_reset_n),
      .col_s1_write_n                                              (col_s1_write_n),
      .col_s1_writedata                                            (col_s1_writedata),
      .cpu_0_data_master_address_to_slave                          (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_col_s1                            (cpu_0_data_master_granted_col_s1),
      .cpu_0_data_master_latency_counter                           (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_col_s1                  (cpu_0_data_master_qualified_request_col_s1),
      .cpu_0_data_master_read                                      (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_col_s1                    (cpu_0_data_master_read_data_valid_col_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_col_s1                           (cpu_0_data_master_requests_col_s1),
      .cpu_0_data_master_write                                     (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                 (cpu_0_data_master_writedata),
      .d1_col_s1_end_xfer                                          (d1_col_s1_end_xfer),
      .reset_n                                                     (clk_0_reset_n)
    );

  col the_col
    (
      .address    (col_s1_address),
      .chipselect (col_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_col),
      .readdata   (col_s1_readdata),
      .reset_n    (col_s1_reset_n),
      .write_n    (col_s1_write_n),
      .writedata  (col_s1_writedata)
    );

  cpu_0_jtag_debug_module_arbitrator the_cpu_0_jtag_debug_module
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                       (cpu_0_data_master_byteenable),
      .cpu_0_data_master_debugaccess                                      (cpu_0_data_master_debugaccess),
      .cpu_0_data_master_granted_cpu_0_jtag_debug_module                  (cpu_0_data_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module        (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module          (cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_cpu_0_jtag_debug_module                 (cpu_0_data_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_cpu_0_jtag_debug_module           (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module   (cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_requests_cpu_0_jtag_debug_module          (cpu_0_instruction_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_jtag_debug_module_address                                    (cpu_0_jtag_debug_module_address),
      .cpu_0_jtag_debug_module_begintransfer                              (cpu_0_jtag_debug_module_begintransfer),
      .cpu_0_jtag_debug_module_byteenable                                 (cpu_0_jtag_debug_module_byteenable),
      .cpu_0_jtag_debug_module_chipselect                                 (cpu_0_jtag_debug_module_chipselect),
      .cpu_0_jtag_debug_module_debugaccess                                (cpu_0_jtag_debug_module_debugaccess),
      .cpu_0_jtag_debug_module_readdata                                   (cpu_0_jtag_debug_module_readdata),
      .cpu_0_jtag_debug_module_readdata_from_sa                           (cpu_0_jtag_debug_module_readdata_from_sa),
      .cpu_0_jtag_debug_module_reset                                      (cpu_0_jtag_debug_module_reset),
      .cpu_0_jtag_debug_module_reset_n                                    (cpu_0_jtag_debug_module_reset_n),
      .cpu_0_jtag_debug_module_resetrequest                               (cpu_0_jtag_debug_module_resetrequest),
      .cpu_0_jtag_debug_module_resetrequest_from_sa                       (cpu_0_jtag_debug_module_resetrequest_from_sa),
      .cpu_0_jtag_debug_module_write                                      (cpu_0_jtag_debug_module_write),
      .cpu_0_jtag_debug_module_writedata                                  (cpu_0_jtag_debug_module_writedata),
      .d1_cpu_0_jtag_debug_module_end_xfer                                (d1_cpu_0_jtag_debug_module_end_xfer),
      .reset_n                                                            (clk_0_reset_n)
    );

  cpu_0_data_master_arbitrator the_cpu_0_data_master
    (
      .button_pio_s1_irq_from_sa                                         (button_pio_s1_irq_from_sa),
      .button_pio_s1_readdata_from_sa                                    (button_pio_s1_readdata_from_sa),
      .cfi_flash_0_s1_wait_counter_eq_0                                  (cfi_flash_0_s1_wait_counter_eq_0),
      .clk                                                               (clk_0),
      .col_s1_readdata_from_sa                                           (col_s1_readdata_from_sa),
      .cpu_0_data_master_address                                         (cpu_0_data_master_address),
      .cpu_0_data_master_address_to_slave                                (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                      (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_cfi_flash_0_s1                       (cpu_0_data_master_byteenable_cfi_flash_0_s1),
      .cpu_0_data_master_byteenable_sdram_0_s1                           (cpu_0_data_master_byteenable_sdram_0_s1),
      .cpu_0_data_master_dbs_address                                     (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                    (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_granted_button_pio_s1                           (cpu_0_data_master_granted_button_pio_s1),
      .cpu_0_data_master_granted_cfi_flash_0_s1                          (cpu_0_data_master_granted_cfi_flash_0_s1),
      .cpu_0_data_master_granted_col_s1                                  (cpu_0_data_master_granted_col_s1),
      .cpu_0_data_master_granted_cpu_0_jtag_debug_module                 (cpu_0_data_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave           (cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_granted_led_pio_s1                              (cpu_0_data_master_granted_led_pio_s1),
      .cpu_0_data_master_granted_row_s1                                  (cpu_0_data_master_granted_row_s1),
      .cpu_0_data_master_granted_sdram_0_s1                              (cpu_0_data_master_granted_sdram_0_s1),
      .cpu_0_data_master_granted_tft_lcd_data_s1                         (cpu_0_data_master_granted_tft_lcd_data_s1),
      .cpu_0_data_master_granted_tft_lcd_nrd_s1                          (cpu_0_data_master_granted_tft_lcd_nrd_s1),
      .cpu_0_data_master_granted_tft_lcd_nrst_s1                         (cpu_0_data_master_granted_tft_lcd_nrst_s1),
      .cpu_0_data_master_granted_tft_lcd_nwr_s1                          (cpu_0_data_master_granted_tft_lcd_nwr_s1),
      .cpu_0_data_master_granted_tft_lcd_rs_s1                           (cpu_0_data_master_granted_tft_lcd_rs_s1),
      .cpu_0_data_master_irq                                             (cpu_0_data_master_irq),
      .cpu_0_data_master_latency_counter                                 (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_button_pio_s1                 (cpu_0_data_master_qualified_request_button_pio_s1),
      .cpu_0_data_master_qualified_request_cfi_flash_0_s1                (cpu_0_data_master_qualified_request_cfi_flash_0_s1),
      .cpu_0_data_master_qualified_request_col_s1                        (cpu_0_data_master_qualified_request_col_s1),
      .cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module       (cpu_0_data_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_qualified_request_led_pio_s1                    (cpu_0_data_master_qualified_request_led_pio_s1),
      .cpu_0_data_master_qualified_request_row_s1                        (cpu_0_data_master_qualified_request_row_s1),
      .cpu_0_data_master_qualified_request_sdram_0_s1                    (cpu_0_data_master_qualified_request_sdram_0_s1),
      .cpu_0_data_master_qualified_request_tft_lcd_data_s1               (cpu_0_data_master_qualified_request_tft_lcd_data_s1),
      .cpu_0_data_master_qualified_request_tft_lcd_nrd_s1                (cpu_0_data_master_qualified_request_tft_lcd_nrd_s1),
      .cpu_0_data_master_qualified_request_tft_lcd_nrst_s1               (cpu_0_data_master_qualified_request_tft_lcd_nrst_s1),
      .cpu_0_data_master_qualified_request_tft_lcd_nwr_s1                (cpu_0_data_master_qualified_request_tft_lcd_nwr_s1),
      .cpu_0_data_master_qualified_request_tft_lcd_rs_s1                 (cpu_0_data_master_qualified_request_tft_lcd_rs_s1),
      .cpu_0_data_master_read                                            (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_button_pio_s1                   (cpu_0_data_master_read_data_valid_button_pio_s1),
      .cpu_0_data_master_read_data_valid_cfi_flash_0_s1                  (cpu_0_data_master_read_data_valid_cfi_flash_0_s1),
      .cpu_0_data_master_read_data_valid_col_s1                          (cpu_0_data_master_read_data_valid_col_s1),
      .cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module         (cpu_0_data_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave   (cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read_data_valid_led_pio_s1                      (cpu_0_data_master_read_data_valid_led_pio_s1),
      .cpu_0_data_master_read_data_valid_row_s1                          (cpu_0_data_master_read_data_valid_row_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1                      (cpu_0_data_master_read_data_valid_sdram_0_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register       (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_data_s1                 (cpu_0_data_master_read_data_valid_tft_lcd_data_s1),
      .cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1                  (cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1),
      .cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1                 (cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1),
      .cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1                  (cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1),
      .cpu_0_data_master_read_data_valid_tft_lcd_rs_s1                   (cpu_0_data_master_read_data_valid_tft_lcd_rs_s1),
      .cpu_0_data_master_readdata                                        (cpu_0_data_master_readdata),
      .cpu_0_data_master_readdatavalid                                   (cpu_0_data_master_readdatavalid),
      .cpu_0_data_master_requests_button_pio_s1                          (cpu_0_data_master_requests_button_pio_s1),
      .cpu_0_data_master_requests_cfi_flash_0_s1                         (cpu_0_data_master_requests_cfi_flash_0_s1),
      .cpu_0_data_master_requests_col_s1                                 (cpu_0_data_master_requests_col_s1),
      .cpu_0_data_master_requests_cpu_0_jtag_debug_module                (cpu_0_data_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave          (cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_requests_led_pio_s1                             (cpu_0_data_master_requests_led_pio_s1),
      .cpu_0_data_master_requests_row_s1                                 (cpu_0_data_master_requests_row_s1),
      .cpu_0_data_master_requests_sdram_0_s1                             (cpu_0_data_master_requests_sdram_0_s1),
      .cpu_0_data_master_requests_tft_lcd_data_s1                        (cpu_0_data_master_requests_tft_lcd_data_s1),
      .cpu_0_data_master_requests_tft_lcd_nrd_s1                         (cpu_0_data_master_requests_tft_lcd_nrd_s1),
      .cpu_0_data_master_requests_tft_lcd_nrst_s1                        (cpu_0_data_master_requests_tft_lcd_nrst_s1),
      .cpu_0_data_master_requests_tft_lcd_nwr_s1                         (cpu_0_data_master_requests_tft_lcd_nwr_s1),
      .cpu_0_data_master_requests_tft_lcd_rs_s1                          (cpu_0_data_master_requests_tft_lcd_rs_s1),
      .cpu_0_data_master_waitrequest                                     (cpu_0_data_master_waitrequest),
      .cpu_0_data_master_write                                           (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                       (cpu_0_data_master_writedata),
      .cpu_0_jtag_debug_module_readdata_from_sa                          (cpu_0_jtag_debug_module_readdata_from_sa),
      .d1_button_pio_s1_end_xfer                                         (d1_button_pio_s1_end_xfer),
      .d1_col_s1_end_xfer                                                (d1_col_s1_end_xfer),
      .d1_cpu_0_jtag_debug_module_end_xfer                               (d1_cpu_0_jtag_debug_module_end_xfer),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                         (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .d1_led_pio_s1_end_xfer                                            (d1_led_pio_s1_end_xfer),
      .d1_row_s1_end_xfer                                                (d1_row_s1_end_xfer),
      .d1_sdram_0_s1_end_xfer                                            (d1_sdram_0_s1_end_xfer),
      .d1_tft_lcd_data_s1_end_xfer                                       (d1_tft_lcd_data_s1_end_xfer),
      .d1_tft_lcd_nrd_s1_end_xfer                                        (d1_tft_lcd_nrd_s1_end_xfer),
      .d1_tft_lcd_nrst_s1_end_xfer                                       (d1_tft_lcd_nrst_s1_end_xfer),
      .d1_tft_lcd_nwr_s1_end_xfer                                        (d1_tft_lcd_nwr_s1_end_xfer),
      .d1_tft_lcd_rs_s1_end_xfer                                         (d1_tft_lcd_rs_s1_end_xfer),
      .d1_tri_state_bridge_0_avalon_slave_end_xfer                       (d1_tri_state_bridge_0_avalon_slave_end_xfer),
      .incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0  (incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                         (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                    (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                 (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .led_pio_s1_readdata_from_sa                                       (led_pio_s1_readdata_from_sa),
      .reset_n                                                           (clk_0_reset_n),
      .row_s1_readdata_from_sa                                           (row_s1_readdata_from_sa),
      .sdram_0_s1_readdata_from_sa                                       (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                    (sdram_0_s1_waitrequest_from_sa),
      .tft_lcd_data_s1_readdata_from_sa                                  (tft_lcd_data_s1_readdata_from_sa),
      .tft_lcd_nrd_s1_readdata_from_sa                                   (tft_lcd_nrd_s1_readdata_from_sa),
      .tft_lcd_nrst_s1_readdata_from_sa                                  (tft_lcd_nrst_s1_readdata_from_sa),
      .tft_lcd_nwr_s1_readdata_from_sa                                   (tft_lcd_nwr_s1_readdata_from_sa),
      .tft_lcd_rs_s1_readdata_from_sa                                    (tft_lcd_rs_s1_readdata_from_sa)
    );

  cpu_0_instruction_master_arbitrator the_cpu_0_instruction_master
    (
      .cfi_flash_0_s1_wait_counter_eq_0                                   (cfi_flash_0_s1_wait_counter_eq_0),
      .clk                                                                (clk_0),
      .cpu_0_instruction_master_address                                   (cpu_0_instruction_master_address),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_dbs_address                               (cpu_0_instruction_master_dbs_address),
      .cpu_0_instruction_master_granted_cfi_flash_0_s1                    (cpu_0_instruction_master_granted_cfi_flash_0_s1),
      .cpu_0_instruction_master_granted_cpu_0_jtag_debug_module           (cpu_0_instruction_master_granted_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_granted_sdram_0_s1                        (cpu_0_instruction_master_granted_sdram_0_s1),
      .cpu_0_instruction_master_granted_tft_lcd_data_s1                   (cpu_0_instruction_master_granted_tft_lcd_data_s1),
      .cpu_0_instruction_master_granted_tft_lcd_nrd_s1                    (cpu_0_instruction_master_granted_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_granted_tft_lcd_nrst_s1                   (cpu_0_instruction_master_granted_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_granted_tft_lcd_nwr_s1                    (cpu_0_instruction_master_granted_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_granted_tft_lcd_rs_s1                     (cpu_0_instruction_master_granted_tft_lcd_rs_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_cfi_flash_0_s1          (cpu_0_instruction_master_qualified_request_cfi_flash_0_s1),
      .cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module (cpu_0_instruction_master_qualified_request_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_qualified_request_sdram_0_s1              (cpu_0_instruction_master_qualified_request_sdram_0_s1),
      .cpu_0_instruction_master_qualified_request_tft_lcd_data_s1         (cpu_0_instruction_master_qualified_request_tft_lcd_data_s1),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1          (cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1         (cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1          (cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1           (cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1            (cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1),
      .cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module   (cpu_0_instruction_master_read_data_valid_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1                (cpu_0_instruction_master_read_data_valid_sdram_0_s1),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1           (cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1            (cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1           (cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1            (cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1             (cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1),
      .cpu_0_instruction_master_readdata                                  (cpu_0_instruction_master_readdata),
      .cpu_0_instruction_master_readdatavalid                             (cpu_0_instruction_master_readdatavalid),
      .cpu_0_instruction_master_requests_cfi_flash_0_s1                   (cpu_0_instruction_master_requests_cfi_flash_0_s1),
      .cpu_0_instruction_master_requests_cpu_0_jtag_debug_module          (cpu_0_instruction_master_requests_cpu_0_jtag_debug_module),
      .cpu_0_instruction_master_requests_sdram_0_s1                       (cpu_0_instruction_master_requests_sdram_0_s1),
      .cpu_0_instruction_master_requests_tft_lcd_data_s1                  (cpu_0_instruction_master_requests_tft_lcd_data_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nrd_s1                   (cpu_0_instruction_master_requests_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nrst_s1                  (cpu_0_instruction_master_requests_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nwr_s1                   (cpu_0_instruction_master_requests_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_requests_tft_lcd_rs_s1                    (cpu_0_instruction_master_requests_tft_lcd_rs_s1),
      .cpu_0_instruction_master_waitrequest                               (cpu_0_instruction_master_waitrequest),
      .cpu_0_jtag_debug_module_readdata_from_sa                           (cpu_0_jtag_debug_module_readdata_from_sa),
      .d1_cpu_0_jtag_debug_module_end_xfer                                (d1_cpu_0_jtag_debug_module_end_xfer),
      .d1_sdram_0_s1_end_xfer                                             (d1_sdram_0_s1_end_xfer),
      .d1_tft_lcd_data_s1_end_xfer                                        (d1_tft_lcd_data_s1_end_xfer),
      .d1_tft_lcd_nrd_s1_end_xfer                                         (d1_tft_lcd_nrd_s1_end_xfer),
      .d1_tft_lcd_nrst_s1_end_xfer                                        (d1_tft_lcd_nrst_s1_end_xfer),
      .d1_tft_lcd_nwr_s1_end_xfer                                         (d1_tft_lcd_nwr_s1_end_xfer),
      .d1_tft_lcd_rs_s1_end_xfer                                          (d1_tft_lcd_rs_s1_end_xfer),
      .d1_tri_state_bridge_0_avalon_slave_end_xfer                        (d1_tri_state_bridge_0_avalon_slave_end_xfer),
      .incoming_data_to_and_from_the_cfi_flash_0                          (incoming_data_to_and_from_the_cfi_flash_0),
      .reset_n                                                            (clk_0_reset_n),
      .sdram_0_s1_readdata_from_sa                                        (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_waitrequest_from_sa                                     (sdram_0_s1_waitrequest_from_sa),
      .tft_lcd_data_s1_readdata_from_sa                                   (tft_lcd_data_s1_readdata_from_sa),
      .tft_lcd_nrd_s1_readdata_from_sa                                    (tft_lcd_nrd_s1_readdata_from_sa),
      .tft_lcd_nrst_s1_readdata_from_sa                                   (tft_lcd_nrst_s1_readdata_from_sa),
      .tft_lcd_nwr_s1_readdata_from_sa                                    (tft_lcd_nwr_s1_readdata_from_sa),
      .tft_lcd_rs_s1_readdata_from_sa                                     (tft_lcd_rs_s1_readdata_from_sa)
    );

  cpu_0 the_cpu_0
    (
      .clk                                   (clk_0),
      .d_address                             (cpu_0_data_master_address),
      .d_byteenable                          (cpu_0_data_master_byteenable),
      .d_irq                                 (cpu_0_data_master_irq),
      .d_read                                (cpu_0_data_master_read),
      .d_readdata                            (cpu_0_data_master_readdata),
      .d_readdatavalid                       (cpu_0_data_master_readdatavalid),
      .d_waitrequest                         (cpu_0_data_master_waitrequest),
      .d_write                               (cpu_0_data_master_write),
      .d_writedata                           (cpu_0_data_master_writedata),
      .i_address                             (cpu_0_instruction_master_address),
      .i_read                                (cpu_0_instruction_master_read),
      .i_readdata                            (cpu_0_instruction_master_readdata),
      .i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),
      .i_waitrequest                         (cpu_0_instruction_master_waitrequest),
      .jtag_debug_module_address             (cpu_0_jtag_debug_module_address),
      .jtag_debug_module_begintransfer       (cpu_0_jtag_debug_module_begintransfer),
      .jtag_debug_module_byteenable          (cpu_0_jtag_debug_module_byteenable),
      .jtag_debug_module_clk                 (clk_0),
      .jtag_debug_module_debugaccess         (cpu_0_jtag_debug_module_debugaccess),
      .jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),
      .jtag_debug_module_readdata            (cpu_0_jtag_debug_module_readdata),
      .jtag_debug_module_reset               (cpu_0_jtag_debug_module_reset),
      .jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_resetrequest),
      .jtag_debug_module_select              (cpu_0_jtag_debug_module_chipselect),
      .jtag_debug_module_write               (cpu_0_jtag_debug_module_write),
      .jtag_debug_module_writedata           (cpu_0_jtag_debug_module_writedata),
      .reset_n                               (cpu_0_jtag_debug_module_reset_n)
    );

  jtag_uart_0_avalon_jtag_slave_arbitrator the_jtag_uart_0_avalon_jtag_slave
    (
      .clk                                                               (clk_0),
      .cpu_0_data_master_address_to_slave                                (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave           (cpu_0_data_master_granted_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_latency_counter                                 (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave (cpu_0_data_master_qualified_request_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read                                            (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave   (cpu_0_data_master_read_data_valid_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register       (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave          (cpu_0_data_master_requests_jtag_uart_0_avalon_jtag_slave),
      .cpu_0_data_master_write                                           (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                       (cpu_0_data_master_writedata),
      .d1_jtag_uart_0_avalon_jtag_slave_end_xfer                         (d1_jtag_uart_0_avalon_jtag_slave_end_xfer),
      .jtag_uart_0_avalon_jtag_slave_address                             (jtag_uart_0_avalon_jtag_slave_address),
      .jtag_uart_0_avalon_jtag_slave_chipselect                          (jtag_uart_0_avalon_jtag_slave_chipselect),
      .jtag_uart_0_avalon_jtag_slave_dataavailable                       (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa               (jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa),
      .jtag_uart_0_avalon_jtag_slave_irq                                 (jtag_uart_0_avalon_jtag_slave_irq),
      .jtag_uart_0_avalon_jtag_slave_irq_from_sa                         (jtag_uart_0_avalon_jtag_slave_irq_from_sa),
      .jtag_uart_0_avalon_jtag_slave_read_n                              (jtag_uart_0_avalon_jtag_slave_read_n),
      .jtag_uart_0_avalon_jtag_slave_readdata                            (jtag_uart_0_avalon_jtag_slave_readdata),
      .jtag_uart_0_avalon_jtag_slave_readdata_from_sa                    (jtag_uart_0_avalon_jtag_slave_readdata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_readyfordata                        (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa                (jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa),
      .jtag_uart_0_avalon_jtag_slave_reset_n                             (jtag_uart_0_avalon_jtag_slave_reset_n),
      .jtag_uart_0_avalon_jtag_slave_waitrequest                         (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa                 (jtag_uart_0_avalon_jtag_slave_waitrequest_from_sa),
      .jtag_uart_0_avalon_jtag_slave_write_n                             (jtag_uart_0_avalon_jtag_slave_write_n),
      .jtag_uart_0_avalon_jtag_slave_writedata                           (jtag_uart_0_avalon_jtag_slave_writedata),
      .reset_n                                                           (clk_0_reset_n)
    );

  jtag_uart_0 the_jtag_uart_0
    (
      .av_address     (jtag_uart_0_avalon_jtag_slave_address),
      .av_chipselect  (jtag_uart_0_avalon_jtag_slave_chipselect),
      .av_irq         (jtag_uart_0_avalon_jtag_slave_irq),
      .av_read_n      (jtag_uart_0_avalon_jtag_slave_read_n),
      .av_readdata    (jtag_uart_0_avalon_jtag_slave_readdata),
      .av_waitrequest (jtag_uart_0_avalon_jtag_slave_waitrequest),
      .av_write_n     (jtag_uart_0_avalon_jtag_slave_write_n),
      .av_writedata   (jtag_uart_0_avalon_jtag_slave_writedata),
      .clk            (clk_0),
      .dataavailable  (jtag_uart_0_avalon_jtag_slave_dataavailable),
      .readyfordata   (jtag_uart_0_avalon_jtag_slave_readyfordata),
      .rst_n          (jtag_uart_0_avalon_jtag_slave_reset_n)
    );

  led_pio_s1_arbitrator the_led_pio_s1
    (
      .clk                                                         (clk_0),
      .cpu_0_data_master_address_to_slave                          (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_led_pio_s1                        (cpu_0_data_master_granted_led_pio_s1),
      .cpu_0_data_master_latency_counter                           (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_led_pio_s1              (cpu_0_data_master_qualified_request_led_pio_s1),
      .cpu_0_data_master_read                                      (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_led_pio_s1                (cpu_0_data_master_read_data_valid_led_pio_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_led_pio_s1                       (cpu_0_data_master_requests_led_pio_s1),
      .cpu_0_data_master_write                                     (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                 (cpu_0_data_master_writedata),
      .d1_led_pio_s1_end_xfer                                      (d1_led_pio_s1_end_xfer),
      .led_pio_s1_address                                          (led_pio_s1_address),
      .led_pio_s1_chipselect                                       (led_pio_s1_chipselect),
      .led_pio_s1_readdata                                         (led_pio_s1_readdata),
      .led_pio_s1_readdata_from_sa                                 (led_pio_s1_readdata_from_sa),
      .led_pio_s1_reset_n                                          (led_pio_s1_reset_n),
      .led_pio_s1_write_n                                          (led_pio_s1_write_n),
      .led_pio_s1_writedata                                        (led_pio_s1_writedata),
      .reset_n                                                     (clk_0_reset_n)
    );

  led_pio the_led_pio
    (
      .address    (led_pio_s1_address),
      .chipselect (led_pio_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_led_pio),
      .readdata   (led_pio_s1_readdata),
      .reset_n    (led_pio_s1_reset_n),
      .write_n    (led_pio_s1_write_n),
      .writedata  (led_pio_s1_writedata)
    );

  row_s1_arbitrator the_row_s1
    (
      .clk                                                         (clk_0),
      .cpu_0_data_master_address_to_slave                          (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_row_s1                            (cpu_0_data_master_granted_row_s1),
      .cpu_0_data_master_latency_counter                           (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_row_s1                  (cpu_0_data_master_qualified_request_row_s1),
      .cpu_0_data_master_read                                      (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_row_s1                    (cpu_0_data_master_read_data_valid_row_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_row_s1                           (cpu_0_data_master_requests_row_s1),
      .cpu_0_data_master_write                                     (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                 (cpu_0_data_master_writedata),
      .d1_row_s1_end_xfer                                          (d1_row_s1_end_xfer),
      .reset_n                                                     (clk_0_reset_n),
      .row_s1_address                                              (row_s1_address),
      .row_s1_chipselect                                           (row_s1_chipselect),
      .row_s1_readdata                                             (row_s1_readdata),
      .row_s1_readdata_from_sa                                     (row_s1_readdata_from_sa),
      .row_s1_reset_n                                              (row_s1_reset_n),
      .row_s1_write_n                                              (row_s1_write_n),
      .row_s1_writedata                                            (row_s1_writedata)
    );

  row the_row
    (
      .address    (row_s1_address),
      .chipselect (row_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_row),
      .readdata   (row_s1_readdata),
      .reset_n    (row_s1_reset_n),
      .write_n    (row_s1_write_n),
      .writedata  (row_s1_writedata)
    );

  sdram_0_s1_arbitrator the_sdram_0_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                       (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_sdram_0_s1                            (cpu_0_data_master_byteenable_sdram_0_s1),
      .cpu_0_data_master_dbs_address                                      (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                     (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_granted_sdram_0_s1                               (cpu_0_data_master_granted_sdram_0_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_sdram_0_s1                     (cpu_0_data_master_qualified_request_sdram_0_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1                       (cpu_0_data_master_read_data_valid_sdram_0_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_sdram_0_s1                              (cpu_0_data_master_requests_sdram_0_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_dbs_address                               (cpu_0_instruction_master_dbs_address),
      .cpu_0_instruction_master_granted_sdram_0_s1                        (cpu_0_instruction_master_granted_sdram_0_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_sdram_0_s1              (cpu_0_instruction_master_qualified_request_sdram_0_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1                (cpu_0_instruction_master_read_data_valid_sdram_0_s1),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_requests_sdram_0_s1                       (cpu_0_instruction_master_requests_sdram_0_s1),
      .d1_sdram_0_s1_end_xfer                                             (d1_sdram_0_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .sdram_0_s1_address                                                 (sdram_0_s1_address),
      .sdram_0_s1_byteenable_n                                            (sdram_0_s1_byteenable_n),
      .sdram_0_s1_chipselect                                              (sdram_0_s1_chipselect),
      .sdram_0_s1_read_n                                                  (sdram_0_s1_read_n),
      .sdram_0_s1_readdata                                                (sdram_0_s1_readdata),
      .sdram_0_s1_readdata_from_sa                                        (sdram_0_s1_readdata_from_sa),
      .sdram_0_s1_readdatavalid                                           (sdram_0_s1_readdatavalid),
      .sdram_0_s1_reset_n                                                 (sdram_0_s1_reset_n),
      .sdram_0_s1_waitrequest                                             (sdram_0_s1_waitrequest),
      .sdram_0_s1_waitrequest_from_sa                                     (sdram_0_s1_waitrequest_from_sa),
      .sdram_0_s1_write_n                                                 (sdram_0_s1_write_n),
      .sdram_0_s1_writedata                                               (sdram_0_s1_writedata)
    );

  sdram_0 the_sdram_0
    (
      .az_addr        (sdram_0_s1_address),
      .az_be_n        (sdram_0_s1_byteenable_n),
      .az_cs          (sdram_0_s1_chipselect),
      .az_data        (sdram_0_s1_writedata),
      .az_rd_n        (sdram_0_s1_read_n),
      .az_wr_n        (sdram_0_s1_write_n),
      .clk            (clk_0),
      .reset_n        (sdram_0_s1_reset_n),
      .za_data        (sdram_0_s1_readdata),
      .za_valid       (sdram_0_s1_readdatavalid),
      .za_waitrequest (sdram_0_s1_waitrequest),
      .zs_addr        (zs_addr_from_the_sdram_0),
      .zs_ba          (zs_ba_from_the_sdram_0),
      .zs_cas_n       (zs_cas_n_from_the_sdram_0),
      .zs_cke         (zs_cke_from_the_sdram_0),
      .zs_cs_n        (zs_cs_n_from_the_sdram_0),
      .zs_dq          (zs_dq_to_and_from_the_sdram_0),
      .zs_dqm         (zs_dqm_from_the_sdram_0),
      .zs_ras_n       (zs_ras_n_from_the_sdram_0),
      .zs_we_n        (zs_we_n_from_the_sdram_0)
    );

  tft_lcd_data_s1_arbitrator the_tft_lcd_data_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                       (cpu_0_data_master_byteenable),
      .cpu_0_data_master_granted_tft_lcd_data_s1                          (cpu_0_data_master_granted_tft_lcd_data_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_tft_lcd_data_s1                (cpu_0_data_master_qualified_request_tft_lcd_data_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_data_s1                  (cpu_0_data_master_read_data_valid_tft_lcd_data_s1),
      .cpu_0_data_master_requests_tft_lcd_data_s1                         (cpu_0_data_master_requests_tft_lcd_data_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_tft_lcd_data_s1                   (cpu_0_instruction_master_granted_tft_lcd_data_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_tft_lcd_data_s1         (cpu_0_instruction_master_qualified_request_tft_lcd_data_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1           (cpu_0_instruction_master_read_data_valid_tft_lcd_data_s1),
      .cpu_0_instruction_master_requests_tft_lcd_data_s1                  (cpu_0_instruction_master_requests_tft_lcd_data_s1),
      .d1_tft_lcd_data_s1_end_xfer                                        (d1_tft_lcd_data_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .tft_lcd_data_s1_address                                            (tft_lcd_data_s1_address),
      .tft_lcd_data_s1_chipselect                                         (tft_lcd_data_s1_chipselect),
      .tft_lcd_data_s1_readdata                                           (tft_lcd_data_s1_readdata),
      .tft_lcd_data_s1_readdata_from_sa                                   (tft_lcd_data_s1_readdata_from_sa),
      .tft_lcd_data_s1_reset_n                                            (tft_lcd_data_s1_reset_n),
      .tft_lcd_data_s1_write_n                                            (tft_lcd_data_s1_write_n),
      .tft_lcd_data_s1_writedata                                          (tft_lcd_data_s1_writedata)
    );

  tft_lcd_data the_tft_lcd_data
    (
      .address    (tft_lcd_data_s1_address),
      .chipselect (tft_lcd_data_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_tft_lcd_data),
      .readdata   (tft_lcd_data_s1_readdata),
      .reset_n    (tft_lcd_data_s1_reset_n),
      .write_n    (tft_lcd_data_s1_write_n),
      .writedata  (tft_lcd_data_s1_writedata)
    );

  tft_lcd_nrd_s1_arbitrator the_tft_lcd_nrd_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_tft_lcd_nrd_s1                           (cpu_0_data_master_granted_tft_lcd_nrd_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_tft_lcd_nrd_s1                 (cpu_0_data_master_qualified_request_tft_lcd_nrd_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1                   (cpu_0_data_master_read_data_valid_tft_lcd_nrd_s1),
      .cpu_0_data_master_requests_tft_lcd_nrd_s1                          (cpu_0_data_master_requests_tft_lcd_nrd_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_tft_lcd_nrd_s1                    (cpu_0_instruction_master_granted_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1          (cpu_0_instruction_master_qualified_request_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1            (cpu_0_instruction_master_read_data_valid_tft_lcd_nrd_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nrd_s1                   (cpu_0_instruction_master_requests_tft_lcd_nrd_s1),
      .d1_tft_lcd_nrd_s1_end_xfer                                         (d1_tft_lcd_nrd_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .tft_lcd_nrd_s1_address                                             (tft_lcd_nrd_s1_address),
      .tft_lcd_nrd_s1_chipselect                                          (tft_lcd_nrd_s1_chipselect),
      .tft_lcd_nrd_s1_readdata                                            (tft_lcd_nrd_s1_readdata),
      .tft_lcd_nrd_s1_readdata_from_sa                                    (tft_lcd_nrd_s1_readdata_from_sa),
      .tft_lcd_nrd_s1_reset_n                                             (tft_lcd_nrd_s1_reset_n),
      .tft_lcd_nrd_s1_write_n                                             (tft_lcd_nrd_s1_write_n),
      .tft_lcd_nrd_s1_writedata                                           (tft_lcd_nrd_s1_writedata)
    );

  tft_lcd_nrd the_tft_lcd_nrd
    (
      .address    (tft_lcd_nrd_s1_address),
      .chipselect (tft_lcd_nrd_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_tft_lcd_nrd),
      .readdata   (tft_lcd_nrd_s1_readdata),
      .reset_n    (tft_lcd_nrd_s1_reset_n),
      .write_n    (tft_lcd_nrd_s1_write_n),
      .writedata  (tft_lcd_nrd_s1_writedata)
    );

  tft_lcd_nrst_s1_arbitrator the_tft_lcd_nrst_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_tft_lcd_nrst_s1                          (cpu_0_data_master_granted_tft_lcd_nrst_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_tft_lcd_nrst_s1                (cpu_0_data_master_qualified_request_tft_lcd_nrst_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1                  (cpu_0_data_master_read_data_valid_tft_lcd_nrst_s1),
      .cpu_0_data_master_requests_tft_lcd_nrst_s1                         (cpu_0_data_master_requests_tft_lcd_nrst_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_tft_lcd_nrst_s1                   (cpu_0_instruction_master_granted_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1         (cpu_0_instruction_master_qualified_request_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1           (cpu_0_instruction_master_read_data_valid_tft_lcd_nrst_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nrst_s1                  (cpu_0_instruction_master_requests_tft_lcd_nrst_s1),
      .d1_tft_lcd_nrst_s1_end_xfer                                        (d1_tft_lcd_nrst_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .tft_lcd_nrst_s1_address                                            (tft_lcd_nrst_s1_address),
      .tft_lcd_nrst_s1_chipselect                                         (tft_lcd_nrst_s1_chipselect),
      .tft_lcd_nrst_s1_readdata                                           (tft_lcd_nrst_s1_readdata),
      .tft_lcd_nrst_s1_readdata_from_sa                                   (tft_lcd_nrst_s1_readdata_from_sa),
      .tft_lcd_nrst_s1_reset_n                                            (tft_lcd_nrst_s1_reset_n),
      .tft_lcd_nrst_s1_write_n                                            (tft_lcd_nrst_s1_write_n),
      .tft_lcd_nrst_s1_writedata                                          (tft_lcd_nrst_s1_writedata)
    );

  tft_lcd_nrst the_tft_lcd_nrst
    (
      .address    (tft_lcd_nrst_s1_address),
      .chipselect (tft_lcd_nrst_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_tft_lcd_nrst),
      .readdata   (tft_lcd_nrst_s1_readdata),
      .reset_n    (tft_lcd_nrst_s1_reset_n),
      .write_n    (tft_lcd_nrst_s1_write_n),
      .writedata  (tft_lcd_nrst_s1_writedata)
    );

  tft_lcd_nwr_s1_arbitrator the_tft_lcd_nwr_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_tft_lcd_nwr_s1                           (cpu_0_data_master_granted_tft_lcd_nwr_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_tft_lcd_nwr_s1                 (cpu_0_data_master_qualified_request_tft_lcd_nwr_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1                   (cpu_0_data_master_read_data_valid_tft_lcd_nwr_s1),
      .cpu_0_data_master_requests_tft_lcd_nwr_s1                          (cpu_0_data_master_requests_tft_lcd_nwr_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_tft_lcd_nwr_s1                    (cpu_0_instruction_master_granted_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1          (cpu_0_instruction_master_qualified_request_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1            (cpu_0_instruction_master_read_data_valid_tft_lcd_nwr_s1),
      .cpu_0_instruction_master_requests_tft_lcd_nwr_s1                   (cpu_0_instruction_master_requests_tft_lcd_nwr_s1),
      .d1_tft_lcd_nwr_s1_end_xfer                                         (d1_tft_lcd_nwr_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .tft_lcd_nwr_s1_address                                             (tft_lcd_nwr_s1_address),
      .tft_lcd_nwr_s1_chipselect                                          (tft_lcd_nwr_s1_chipselect),
      .tft_lcd_nwr_s1_readdata                                            (tft_lcd_nwr_s1_readdata),
      .tft_lcd_nwr_s1_readdata_from_sa                                    (tft_lcd_nwr_s1_readdata_from_sa),
      .tft_lcd_nwr_s1_reset_n                                             (tft_lcd_nwr_s1_reset_n),
      .tft_lcd_nwr_s1_write_n                                             (tft_lcd_nwr_s1_write_n),
      .tft_lcd_nwr_s1_writedata                                           (tft_lcd_nwr_s1_writedata)
    );

  tft_lcd_nwr the_tft_lcd_nwr
    (
      .address    (tft_lcd_nwr_s1_address),
      .chipselect (tft_lcd_nwr_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_tft_lcd_nwr),
      .readdata   (tft_lcd_nwr_s1_readdata),
      .reset_n    (tft_lcd_nwr_s1_reset_n),
      .write_n    (tft_lcd_nwr_s1_write_n),
      .writedata  (tft_lcd_nwr_s1_writedata)
    );

  tft_lcd_rs_s1_arbitrator the_tft_lcd_rs_s1
    (
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_granted_tft_lcd_rs_s1                            (cpu_0_data_master_granted_tft_lcd_rs_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_tft_lcd_rs_s1                  (cpu_0_data_master_qualified_request_tft_lcd_rs_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_read_data_valid_tft_lcd_rs_s1                    (cpu_0_data_master_read_data_valid_tft_lcd_rs_s1),
      .cpu_0_data_master_requests_tft_lcd_rs_s1                           (cpu_0_data_master_requests_tft_lcd_rs_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_data_master_writedata                                        (cpu_0_data_master_writedata),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_granted_tft_lcd_rs_s1                     (cpu_0_instruction_master_granted_tft_lcd_rs_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1           (cpu_0_instruction_master_qualified_request_tft_lcd_rs_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1             (cpu_0_instruction_master_read_data_valid_tft_lcd_rs_s1),
      .cpu_0_instruction_master_requests_tft_lcd_rs_s1                    (cpu_0_instruction_master_requests_tft_lcd_rs_s1),
      .d1_tft_lcd_rs_s1_end_xfer                                          (d1_tft_lcd_rs_s1_end_xfer),
      .reset_n                                                            (clk_0_reset_n),
      .tft_lcd_rs_s1_address                                              (tft_lcd_rs_s1_address),
      .tft_lcd_rs_s1_chipselect                                           (tft_lcd_rs_s1_chipselect),
      .tft_lcd_rs_s1_readdata                                             (tft_lcd_rs_s1_readdata),
      .tft_lcd_rs_s1_readdata_from_sa                                     (tft_lcd_rs_s1_readdata_from_sa),
      .tft_lcd_rs_s1_reset_n                                              (tft_lcd_rs_s1_reset_n),
      .tft_lcd_rs_s1_write_n                                              (tft_lcd_rs_s1_write_n),
      .tft_lcd_rs_s1_writedata                                            (tft_lcd_rs_s1_writedata)
    );

  tft_lcd_rs the_tft_lcd_rs
    (
      .address    (tft_lcd_rs_s1_address),
      .chipselect (tft_lcd_rs_s1_chipselect),
      .clk        (clk_0),
      .out_port   (out_port_from_the_tft_lcd_rs),
      .readdata   (tft_lcd_rs_s1_readdata),
      .reset_n    (tft_lcd_rs_s1_reset_n),
      .write_n    (tft_lcd_rs_s1_write_n),
      .writedata  (tft_lcd_rs_s1_writedata)
    );

  tri_state_bridge_0_avalon_slave_arbitrator the_tri_state_bridge_0_avalon_slave
    (
      .address_to_the_cfi_flash_0                                         (address_to_the_cfi_flash_0),
      .cfi_flash_0_s1_wait_counter_eq_0                                   (cfi_flash_0_s1_wait_counter_eq_0),
      .clk                                                                (clk_0),
      .cpu_0_data_master_address_to_slave                                 (cpu_0_data_master_address_to_slave),
      .cpu_0_data_master_byteenable                                       (cpu_0_data_master_byteenable),
      .cpu_0_data_master_byteenable_cfi_flash_0_s1                        (cpu_0_data_master_byteenable_cfi_flash_0_s1),
      .cpu_0_data_master_dbs_address                                      (cpu_0_data_master_dbs_address),
      .cpu_0_data_master_dbs_write_16                                     (cpu_0_data_master_dbs_write_16),
      .cpu_0_data_master_granted_cfi_flash_0_s1                           (cpu_0_data_master_granted_cfi_flash_0_s1),
      .cpu_0_data_master_latency_counter                                  (cpu_0_data_master_latency_counter),
      .cpu_0_data_master_qualified_request_cfi_flash_0_s1                 (cpu_0_data_master_qualified_request_cfi_flash_0_s1),
      .cpu_0_data_master_read                                             (cpu_0_data_master_read),
      .cpu_0_data_master_read_data_valid_cfi_flash_0_s1                   (cpu_0_data_master_read_data_valid_cfi_flash_0_s1),
      .cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register        (cpu_0_data_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_data_master_requests_cfi_flash_0_s1                          (cpu_0_data_master_requests_cfi_flash_0_s1),
      .cpu_0_data_master_write                                            (cpu_0_data_master_write),
      .cpu_0_instruction_master_address_to_slave                          (cpu_0_instruction_master_address_to_slave),
      .cpu_0_instruction_master_dbs_address                               (cpu_0_instruction_master_dbs_address),
      .cpu_0_instruction_master_granted_cfi_flash_0_s1                    (cpu_0_instruction_master_granted_cfi_flash_0_s1),
      .cpu_0_instruction_master_latency_counter                           (cpu_0_instruction_master_latency_counter),
      .cpu_0_instruction_master_qualified_request_cfi_flash_0_s1          (cpu_0_instruction_master_qualified_request_cfi_flash_0_s1),
      .cpu_0_instruction_master_read                                      (cpu_0_instruction_master_read),
      .cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1            (cpu_0_instruction_master_read_data_valid_cfi_flash_0_s1),
      .cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register (cpu_0_instruction_master_read_data_valid_sdram_0_s1_shift_register),
      .cpu_0_instruction_master_requests_cfi_flash_0_s1                   (cpu_0_instruction_master_requests_cfi_flash_0_s1),
      .d1_tri_state_bridge_0_avalon_slave_end_xfer                        (d1_tri_state_bridge_0_avalon_slave_end_xfer),
      .data_to_and_from_the_cfi_flash_0                                   (data_to_and_from_the_cfi_flash_0),
      .incoming_data_to_and_from_the_cfi_flash_0                          (incoming_data_to_and_from_the_cfi_flash_0),
      .incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0   (incoming_data_to_and_from_the_cfi_flash_0_with_Xs_converted_to_0),
      .read_n_to_the_cfi_flash_0                                          (read_n_to_the_cfi_flash_0),
      .reset_n                                                            (clk_0_reset_n),
      .select_n_to_the_cfi_flash_0                                        (select_n_to_the_cfi_flash_0),
      .write_n_to_the_cfi_flash_0                                         (write_n_to_the_cfi_flash_0)
    );

  //reset is asserted asynchronously and deasserted synchronously
  nioscpu_reset_clk_0_domain_synch_module nioscpu_reset_clk_0_domain_synch
    (
      .clk      (clk_0),
      .data_in  (1'b1),
      .data_out (clk_0_reset_n),
      .reset_n  (reset_n_sources)
    );

  //reset sources mux, which is an e_mux
  assign reset_n_sources = ~(~reset_n |
    0 |
    cpu_0_jtag_debug_module_resetrequest_from_sa |
    cpu_0_jtag_debug_module_resetrequest_from_sa);


endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cfi_flash_0_lane0_module (
                                  // inputs:
                                   data,
                                   rdaddress,
                                   rdclken,
                                   wraddress,
                                   wrclock,
                                   wren,

                                  // outputs:
                                   q
                                )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 20: 0] rdaddress;
  input            rdclken;
  input   [ 20: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [2097151: 0];
  wire    [  7: 0] q;
  reg     [ 20: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("cfi_flash_0_lane0.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "cfi_flash_0_lane0.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 21,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cfi_flash_0_lane1_module (
                                  // inputs:
                                   data,
                                   rdaddress,
                                   rdclken,
                                   wraddress,
                                   wrclock,
                                   wren,

                                  // outputs:
                                   q
                                )
;

  output  [  7: 0] q;
  input   [  7: 0] data;
  input   [ 20: 0] rdaddress;
  input            rdclken;
  input   [ 20: 0] wraddress;
  input            wrclock;
  input            wren;

  reg     [  7: 0] mem_array [2097151: 0];
  wire    [  7: 0] q;
  reg     [ 20: 0] read_address;

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  always @(rdaddress)
    begin
      read_address = rdaddress;
    end


  // Data read is asynchronous.
  assign q = mem_array[read_address];

initial
    $readmemh("cfi_flash_0_lane1.dat", mem_array);
  always @(posedge wrclock)
    begin
      // Write data
      if (wren)
          mem_array[wraddress] <= data;
    end



//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on
//synthesis read_comments_as_HDL on
//  always @(rdaddress)
//    begin
//      read_address = rdaddress;
//    end
//
//
//  lpm_ram_dp lpm_ram_dp_component
//    (
//      .data (data),
//      .q (q),
//      .rdaddress (read_address),
//      .rdclken (rdclken),
//      .wraddress (wraddress),
//      .wrclock (wrclock),
//      .wren (wren)
//    );
//
//  defparam lpm_ram_dp_component.lpm_file = "cfi_flash_0_lane1.mif",
//           lpm_ram_dp_component.lpm_hint = "USE_EAB=ON",
//           lpm_ram_dp_component.lpm_indata = "REGISTERED",
//           lpm_ram_dp_component.lpm_outdata = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_rdaddress_control = "UNREGISTERED",
//           lpm_ram_dp_component.lpm_width = 8,
//           lpm_ram_dp_component.lpm_widthad = 21,
//           lpm_ram_dp_component.lpm_wraddress_control = "REGISTERED",
//           lpm_ram_dp_component.suppress_memory_conversion_warnings = "ON";
//
//synthesis read_comments_as_HDL off

endmodule



// turn off superfluous verilog processor warnings 
// altera message_level Level1 
// altera message_off 10034 10035 10036 10037 10230 10240 10030 

module cfi_flash_0 (
                     // inputs:
                      address,
                      read_n,
                      select_n,
                      write_n,

                     // outputs:
                      data
                   )
;

  inout   [ 15: 0] data;
  input   [ 20: 0] address;
  input            read_n;
  input            select_n;
  input            write_n;

  wire    [ 15: 0] data;
  wire    [  7: 0] data_0;
  wire    [  7: 0] data_1;
  wire    [ 15: 0] logic_vector_gasket;
  wire    [  7: 0] q_0;
  wire    [  7: 0] q_1;
  //s1, which is an e_ptf_slave

//synthesis translate_off
//////////////// SIMULATION-ONLY CONTENTS
  assign logic_vector_gasket = data;
  assign data_0 = logic_vector_gasket[7 : 0];
  //cfi_flash_0_lane0, which is an e_ram
  cfi_flash_0_lane0_module cfi_flash_0_lane0
    (
      .data      (data_0),
      .q         (q_0),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data_1 = logic_vector_gasket[15 : 8];
  //cfi_flash_0_lane1, which is an e_ram
  cfi_flash_0_lane1_module cfi_flash_0_lane1
    (
      .data      (data_1),
      .q         (q_1),
      .rdaddress (address),
      .rdclken   (1'b1),
      .wraddress (address),
      .wrclock   (write_n),
      .wren      (~select_n)
    );

  assign data = (~select_n & ~read_n)? {q_1,
    q_0}: {16{1'bz}};


//////////////// END SIMULATION-ONLY CONTENTS

//synthesis translate_on

endmodule


//synthesis translate_off



// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE

// AND HERE WILL BE PRESERVED </ALTERA_NOTE>


// If user logic components use Altsync_Ram with convert_hex2ver.dll,
// set USE_convert_hex2ver in the user comments section above

// `ifdef USE_convert_hex2ver
// `else
// `define NO_PLI 1
// `endif

`include "c:/altera/90/quartus/eda/sim_lib/altera_mf.v"
`include "c:/altera/90/quartus/eda/sim_lib/220model.v"
`include "c:/altera/90/quartus/eda/sim_lib/sgate.v"
`include "sdram_0.v"
`include "sdram_0_test_component.v"
`include "cpu_0_test_bench.v"
`include "cpu_0_mult_cell.v"
`include "cpu_0_oci_test_bench.v"
`include "cpu_0_jtag_debug_module_tck.v"
`include "cpu_0_jtag_debug_module_sysclk.v"
`include "cpu_0_jtag_debug_module_wrapper.v"
`include "cpu_0.v"
`include "button_pio.v"
`include "tft_lcd_nwr.v"
`include "tft_lcd_nrst.v"
`include "tft_lcd_data.v"
`include "row.v"
`include "col.v"
`include "led_pio.v"
`include "jtag_uart_0.v"
`include "tft_lcd_nrd.v"
`include "tft_lcd_rs.v"

`timescale 1ns / 1ps

module test_bench 
;


  wire    [ 21: 0] address_to_the_cfi_flash_0;
  wire             clk;
  reg              clk_0;
  wire    [ 15: 0] data_to_and_from_the_cfi_flash_0;
  wire    [  7: 0] in_port_to_the_button_pio;
  wire             jtag_uart_0_avalon_jtag_slave_dataavailable_from_sa;
  wire             jtag_uart_0_avalon_jtag_slave_readyfordata_from_sa;
  wire    [  3: 0] out_port_from_the_col;
  wire    [  7: 0] out_port_from_the_led_pio;
  wire    [ 15: 0] out_port_from_the_row;
  wire    [  7: 0] out_port_from_the_tft_lcd_data;
  wire             out_port_from_the_tft_lcd_nrd;
  wire             out_port_from_the_tft_lcd_nrst;
  wire             out_port_from_the_tft_lcd_nwr;
  wire             out_port_from_the_tft_lcd_rs;
  wire             read_n_to_the_cfi_flash_0;
  reg              reset_n;
  wire             select_n_to_the_cfi_flash_0;
  wire             write_n_to_the_cfi_flash_0;
  wire    [ 11: 0] zs_addr_from_the_sdram_0;
  wire    [  1: 0] zs_ba_from_the_sdram_0;
  wire             zs_cas_n_from_the_sdram_0;
  wire             zs_cke_from_the_sdram_0;
  wire             zs_cs_n_from_the_sdram_0;
  wire    [ 15: 0] zs_dq_to_and_from_the_sdram_0;
  wire    [  1: 0] zs_dqm_from_the_sdram_0;
  wire             zs_ras_n_from_the_sdram_0;
  wire             zs_we_n_from_the_sdram_0;


// <ALTERA_NOTE> CODE INSERTED BETWEEN HERE
//  add your signals and additional architecture here
// AND HERE WILL BE PRESERVED </ALTERA_NOTE>

  //Set us up the Dut
  nioscpu DUT
    (
      .address_to_the_cfi_flash_0       (address_to_the_cfi_flash_0),
      .clk_0                            (clk_0),
      .data_to_and_from_the_cfi_flash_0 (data_to_and_from_the_cfi_flash_0),
      .in_port_to_the_button_pio        (in_port_to_the_button_pio),
      .out_port_from_the_col            (out_port_from_the_col),
      .out_port_from_the_led_pio        (out_port_from_the_led_pio),
      .out_port_from_the_row            (out_port_from_the_row),
      .out_port_from_the_tft_lcd_data   (out_port_from_the_tft_lcd_data),
      .out_port_from_the_tft_lcd_nrd    (out_port_from_the_tft_lcd_nrd),
      .out_port_from_the_tft_lcd_nrst   (out_port_from_the_tft_lcd_nrst),
      .out_port_from_the_tft_lcd_nwr    (out_port_from_the_tft_lcd_nwr),
      .out_port_from_the_tft_lcd_rs     (out_port_from_the_tft_lcd_rs),
      .read_n_to_the_cfi_flash_0        (read_n_to_the_cfi_flash_0),
      .reset_n                          (reset_n),
      .select_n_to_the_cfi_flash_0      (select_n_to_the_cfi_flash_0),
      .write_n_to_the_cfi_flash_0       (write_n_to_the_cfi_flash_0),
      .zs_addr_from_the_sdram_0         (zs_addr_from_the_sdram_0),
      .zs_ba_from_the_sdram_0           (zs_ba_from_the_sdram_0),
      .zs_cas_n_from_the_sdram_0        (zs_cas_n_from_the_sdram_0),
      .zs_cke_from_the_sdram_0          (zs_cke_from_the_sdram_0),
      .zs_cs_n_from_the_sdram_0         (zs_cs_n_from_the_sdram_0),
      .zs_dq_to_and_from_the_sdram_0    (zs_dq_to_and_from_the_sdram_0),
      .zs_dqm_from_the_sdram_0          (zs_dqm_from_the_sdram_0),
      .zs_ras_n_from_the_sdram_0        (zs_ras_n_from_the_sdram_0),
      .zs_we_n_from_the_sdram_0         (zs_we_n_from_the_sdram_0)
    );

  cfi_flash_0 the_cfi_flash_0
    (
      .address  (address_to_the_cfi_flash_0[21 : 1]),
      .data     (data_to_and_from_the_cfi_flash_0),
      .read_n   (read_n_to_the_cfi_flash_0),
      .select_n (select_n_to_the_cfi_flash_0),
      .write_n  (write_n_to_the_cfi_flash_0)
    );

  sdram_0_test_component the_sdram_0_test_component
    (
      .clk      (clk_0),
      .zs_addr  (zs_addr_from_the_sdram_0),
      .zs_ba    (zs_ba_from_the_sdram_0),
      .zs_cas_n (zs_cas_n_from_the_sdram_0),
      .zs_cke   (zs_cke_from_the_sdram_0),
      .zs_cs_n  (zs_cs_n_from_the_sdram_0),
      .zs_dq    (zs_dq_to_and_from_the_sdram_0),
      .zs_dqm   (zs_dqm_from_the_sdram_0),
      .zs_ras_n (zs_ras_n_from_the_sdram_0),
      .zs_we_n  (zs_we_n_from_the_sdram_0)
    );

  initial
    clk_0 = 1'b0;
  always
    #10 clk_0 <= ~clk_0;
  
  initial 
    begin
      reset_n <= 0;
      #200 reset_n <= 1;
    end

endmodule


//synthesis translate_on