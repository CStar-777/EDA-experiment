module dot_matrix1(clk,reset,row,col);
input clk,reset;
output reg [15:0]row;      //�� 
output reg [3:0]col;       //��
reg [15:0] count1;
reg [31:0] count2;
reg clk_500,divi_1hz;
reg [1:0]cnt4;

always @(posedge clk)
	if(count1==50000000/(5000*2)-1)
		begin
			clk_500 <= ~clk_500;
			count1 <= 16'd0;
		end
	else
		begin
			count1 <= count1 + 16'd1;
		end

always @(posedge clk) begin
	if (count2 == 24999999) begin 
		divi_1hz <= !divi_1hz;
		count2 <= 0;
	end
	else begin
		count2 = count2 + 1;
	end
end

always @(posedge divi_1hz)
	cnt4=cnt4+1;

/***************�ַ���ʾ*******************/ 
initial col=4'b0;
always @(posedge clk_500) begin
	if (!reset)    col<=4'b0;
	else 
	begin      //���ü����������е�  16 �ֱ��룺0000-1111
		if(col==4'b1111) col<=4'b0;
		else col<=col+1;
	end
end

always @(reset or col)begin
	if (!reset)  row<=16'b0; 
	else
	begin 
		if(cnt4 == 2'b00) // xue
		begin
			case (col)
			4'b0000: row <= 16'h7FFF; //�� 1 ��
			4'b0001: row <= 16'h4008; //�� 2 ��
			4'b0010: row <= 16'h4208; //�� 3 ��
			4'b0011: row <= 16'h5D8C; //�� 4 ��
			4'b0100: row <= 16'h6079; //�� 5 ��
			4'b0101: row <= 16'h0082; //�� 6 ��
			4'b0110: row <= 16'h10C4; //�� 7 ��
			4'b0111: row <= 16'h1398; //�� 8 ��
			4'b1000: row <= 16'h0C90; //�� 9 ��
			4'b1001: row <= 16'hF080; //�� 10 ��
			4'b1010: row <= 16'h5080; //�� 11 ��
			4'b1011: row <= 16'h17FF; //�� 12 ��
			4'b1100: row <= 16'h1080; //�� 13 ��
			4'b1101: row <= 16'h1090; //�� 14 ��
			4'b1110: row <= 16'h1088; //�� 15 ��
			4'b1111: row <= 16'h1086; //�� 16 ��
			endcase
		end
		else if(cnt4 == 2'b01) // jie
		begin
			case (col)
			4'b0000: row <= 16'h0010; //�� 1 ��
			4'b0001: row <= 16'h0062; //�� 2 ��
			4'b0010: row <= 16'h47a2; //�� 3 ��
			4'b0011: row <= 16'h5524; //�� 4 ��
			4'b0100: row <= 16'h5564; //�� 5 ��
			4'b0101: row <= 16'hf36f; //�� 6 ��
			4'b0110: row <= 16'h5555; //�� 7 ��
			4'b0111: row <= 16'h5555; //�� 8 ��
			4'b1000: row <= 16'h57fd; //�� 9 ��
			4'b1001: row <= 16'h04e5; //�� 10 ��
			4'b1010: row <= 16'h0d55; //�� 11 ��
			4'b1011: row <= 16'hfb6d; //�� 12 ��
			4'b1100: row <= 16'h8a6f; //�� 13 ��
			4'b1101: row <= 16'h8a64; //�� 14 ��
			4'b1110: row <= 16'hf524; //�� 15 ��
			4'b1111: row <= 16'h1926; //�� 16 ��
			endcase
		end
		else if(cnt4 == 2'b10) // piao
		begin
			case (col)
			4'b0000: row <= 16'h7ff8; //�� 1 ��
			4'b0001: row <= 16'h4020; //�� 2 ��
			4'b0010: row <= 16'h4020; //�� 3 ��
			4'b0011: row <= 16'h7ff0; //�� 4 ��
			4'b0100: row <= 16'h0000; //�� 5 ��
			4'b0101: row <= 16'h8000; //�� 6 ��
			4'b0110: row <= 16'hffff; //�� 7 ��
			4'b0111: row <= 16'h8e18; //�� 8 ��
			4'b1000: row <= 16'hf198; //�� 9 ��
			4'b1001: row <= 16'h4070; //�� 10 ��
			4'b1010: row <= 16'h8ff0; //�� 11 ��
			4'b1011: row <= 16'h8820; //�� 12 ��
			4'b1100: row <= 16'h8820; //�� 13 ��
			4'b1101: row <= 16'h8ff0; //�� 14 ��
			4'b1110: row <= 16'h8000; //�� 15 ��
			4'b1111: row <= 16'h7fff; //�� 16 ��
			endcase
		end
		else if(cnt4 == 2'b11) // liang
		begin
			case (col)
			4'b0000: row <= 16'h0001; //�� 1 ��
			4'b0001: row <= 16'h0202; //�� 2 ��
			4'b0010: row <= 16'hc204; //�� 3 ��
			4'b0011: row <= 16'h63fc; //�� 4 ��
			4'b0100: row <= 16'h0202; //�� 5 ��
			4'b0101: row <= 16'h0002; //�� 6 ��
			4'b0110: row <= 16'h0005; //�� 7 ��
			4'b0111: row <= 16'h1009; //�� 8 ��
			4'b1000: row <= 16'h1209; //�� 9 ��
			4'b1001: row <= 16'h1110; //�� 10 ��
			4'b1010: row <= 16'hd0a0; //�� 11 ��
			4'b1011: row <= 16'h70c0; //�� 12 ��
			4'b1100: row <= 16'h13e0; //�� 13 ��
			4'b1101: row <= 16'h0e30; //�� 14 ��
			4'b1110: row <= 16'h1018; //�� 15 ��
			4'b1111: row <= 16'h100c; //�� 16 ��
			endcase
		end
	end
end
endmodule
 